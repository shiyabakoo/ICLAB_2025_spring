../00_TESTBED/TESTBED.sv