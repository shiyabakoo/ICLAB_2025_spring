`define CYCLE_TIME 11.6

module PATTERN(
    clk,
    rst_n,
    in_valid,
    in_valid2,
    in_data,
    out_valid,
    out_sad
);
output reg clk, rst_n, in_valid, in_valid2;
output reg [11:0] in_data;
input out_valid;
input out_sad;


`protected
b29\GVSSc@>.2KEPOE5aL@6A5BU#^G9#MaMeR#X>7,]g.7J^c/C#/)c+2B?8I;XF
dUfOXE;L.)V#3g_\51:J2&G;3L]QS=+\Ic^B)Y0X.=/A-G[VW_[aOT\]d#D#Z-7d
\-(gg2L]38d,.Af.7<V#2I&7(Y96LefYNVKXSN70;gOM6F.]YS#6\/4F+NbW6C+=
4eC(]FEXDCFX@[+cA+dL;SE/V.CgP,K[]O9ZgO1RRL=fb@fBV5+/5VEXL4c7Jg+O
5b:aW<];AAVa2IbFgTE0#aE:N1/BUK3B5@@<72D\3)9>eX9@EK#=7C_U]5NDc4C?
b+];F76TM)gJ1Ie>GX_;PL;=8BM:OcZg13.>5Ng&DYe9VSS?U;^:b<6BV=+;VB,W
XfMU0\#RH]#\FHb8O8IZg+Q#>XDS0/f>&2(\(g?FJ-OY;]X6?:@2=DO<=\55C2c+
GAC>61MZJcL27c]<\,O\Z0TQ<_3HF:,GgV^<=BfBfJD<&H-dSE^c/,AA9Z3B@4T[
)W=Q7UB?+?UQN[](,P9MCR=U7AcZ/)5H9URNRQ@=e6g\[)[Y2910?a9</CKIK.U,
0&4TEPF:<bgdSe>OMX^0-FPROX@Wa=02=eU3_Wef6e:DSIdW.9^\WIUMH[fN_+W.
/F3c3=7&I_7WaW]9&YM1.@^?^X6K8CUQ+_c/>U^#YIf148XFJdHC0a].Y7U6W)Qc
_@.DPbJ:IR4XF)QXO4#/_->3YK&J0_T#?W,W)VOdXA;fP\N-R/IHd7SGOT>A0eA,
._BD_2XWBS1C\42R6U5_CLS+T0^,_g:TGg7a=[62V-WJ5OZOI?TdF_W,^H/43M6R
4)_;f.#9RX2PT1V8^N#LJLI0GD<K4Z-?g:QI>=]Sb\&O>#Me4MYf#IPNX<B5O9)]
A:f9F94SA:?b3f7Z<@<)L>Zc)R.20>F](E5fTeIE(GWOb3Z27@K@4(Dd0TgBYJJe
NEd6N\aL6)7S4AX?/PD@FS>-bXR.5@1EZ73eB8ZGX/ddgb7:Gcd#9@J:eg@I\Q^U
OSKL?c)5(DL)6VE/A19bT#LbXVI1Y>?)ga/[][-8=2L:;ODg3M,OFNbV/G>7>SAa
K,<BX5a^7fN^]G/XPI9(O>;-@+[7b.KgMWffRBa#<1]IX<a=1P)eM/<.\PXK&IDX
JA/g0M(.O.LE)-\AF>8YWT?.SeH+b@9)^D/V<DTPWSaNBHad+E.:3HIDUHX+)fgP
/9+TLH+/[M8]W.@,7e8<1QAARE^U,9Eb;1:36b5deeXRZeHK2;PPG@FGB.4V3\.b
/3W#-/87:UZE5WLGYMAVX9Mf4[3@7P4g12NFFJ-,;3g-\QfL;W7/2IB4R^+UL]VC
Q\,gAc)0I/Q.U:;HRW)VbNeLDW>[PX.8(0FCg[&dDHIM.3UG/K?fT)9F6A5PaI(J
1N_8FG/@NKZ71[HQ8/eU8@;c3];fBHP.1T?.-7gH664B42I:=5I_gF_/MWM2G6#b
gLRc/4Ha,-&M.7X4Ac5QSL]-U1&[3.HU84NHVcP\gIVB@YJE.AN_N/Y1Wf\>S?6A
fdOEP-L4@;=[^V1ffA2fJC][A-_[M_VTTYS6g-.]URFf8Q.83X(+82cWF.dd&R?S
d<P&&D#E;HE5<7A169E&OYNSIG7W+\[dT6(-aA+=&\K<;HfA4.]+8]0:FZE[P97?
?2N3,d39Z-:3:0?6J;6;^8<Tb9eFJV5SU#S[4cX1W-:Ab2c#F>EQJ#U>98Dd,6I^
Z#=@(gbD,#Q7f[XA/#[HES:@[O;Z&M::<F]#9A1\+)H>0073Y#3^d1PQR+I#fOd]
NKaCVO:LK#/^JL4V_;:U:P_3=+=\__06G#KO803gKgGB-^&Db=?cYM,Mc[G?R8gS
>CD2;0\:(M-=a/-9P0#Hd./TEI>AZYNJ+ceVBVDZ]SQ\M8:OIFbYD-,J3f8;2^IC
2HGDd_/7Eb9;Z9<[,F>,YH]4OA>VG8S[6Ec)?.IQ)Ug94=V(W-cVeDOKX=X,27RR
0e#5[Q?9Z_=<Z)/W[1Q&7\\R(?<I0AM[eBKLI9>Y7OL-bE6BXdI^W>CP<0DcL>>L
Y^.QBHVg_>UfH0^fOO2eV,5fXf8B0WP2\e3_@JS#+Lb:/&CH4621MQ:aL,W.8gg;
7b[7F6YR>O<O>,]0a+g[:A2UEgB41L3)66RY^&;F0PJ9/;G_WGR1EV#+&Jg[O)QG
aA_4P0\H\eg)?:4@6_9dP/)X-@T8>+XXA_VZ]Y#,,KfK)3/X,90OMETZ?b+b#IYS
3#Dd=:U)G4-4K#Q#cRPDEO[81&Z;F;0EV4GE\JfC7B<+HL;(E@Za>D1E.Hd-8;@_
S(4=WX\@Va?O0(6/QXE;fSBJQ53EU8g+)f)Ne<=]UFb5<N6cY<&C8\/D=OIDL4=0
/KN>cY4Z\T;/H#:DB)Q<[I20:d)0\ffaL4U0W^&_&)(#:5A[CK@]]F2;K;d7b8.A
Y05gNBOZ919^UCZKa76B+U::^X[PF8cDKg)++P_F41>ga>G49;498\Y/3SA,R32Y
1,(KK3K)O//b<=HV43J[^g;WA>4UK7AEb.TfM^WNC/)_fUXK5/afe;T3&S7b:L_=
g2+8_&3OFK)_J[IW+46JfHfN5>20Fc@=M5cDO&#Uc=T_cQ=R2-VGQJ8#5Mg0#<+S
&,JeG,EM\:A<,J-+E/->D?g-W\V7_=4IUUQPYDVJSXHK)4XQ&ENCW#B@U#E@IV&W
P11Z?HN0GXQ<48Seb4.QZCAC(O^9&Z=+>:BB=2?>[>3F_GRfS8-7+F]33H6VT^97
#,D:A]:?.4.+OYBO@[DG^#Z11OWDGZ_\e8@XOU>Nd86b=PP._?f9BP\&0#dP6Y8-
7b2NZ&fVE2IXF1/<,6e@O9M+@IPabL;#LDIP]<2Mg&QNIe-HSN=:XAY^c9gIbX6A
(@&A;]aQ_@\0],+Ke[-I2ZGZ&>.BJ1K&</_OS9P_(E&)=2g7<f=KAQKFB:f]c5&H
(.f+<Q5&bgD<I4ZIaBL+N4/We>3TFIcL)NcE/PHX2KNJ;/NcIJVS=8H09\E1&=M[
52PZeCQSReDW/+3=O^d#5G]/Lc[\9a48D#,6@58YGP6^0aACa95H:A1O/OIN7H10
IEPCNPRfYKO=FQ4/LDAF<eAacTbI1-GO>VSOeDM7#f@=6A=U>?aZ.VbW,?SaDEdE
X:EF0GT91<6FS&,?.WQOT-\c/G(74H@4b\PeZgFIFC0/<>gcRf.XDE\;^<cDb(&<
]WZRc5@A5V4=_d7#f55gF?ZB10PF(_#S,K-COT&UC21^7]Z3#5ZA@f7W389BYJ7F
>@PD\4R-fMP(S\D;<B/R_LI)dX6b\MGbD9AVb+A-6N<ROL[_NDW>9<5,A7A-[JX:
be;,I9?R+86P1D\)(0JTcR-MWKf_[T\7;5b;J(H^b(UHTDFNSd(UPeKS5^</I(1S
#B07S683b,^.=V(\EM=V(I,ME3[1/:-MCE+NK+.AbV1]O[^L(^5<:PDQBKfY-d4)
TCQ_9eX;d:L+\gS8W1JR#8+-XJH)@X)<7)/UPMDD:P:SP__f6W]R\OgE</HDZ<LD
#XU-9dCbZCXeXIA&g@ZZQYGeC&NM]IS=UJG<?M@M^edWa5ZW\bD=Bd9QLEW>E,^T
cad&#XF.OdXVZH07UWaMbYg0JQOXd8](A,V^WDcLXJCU(11CO0E7I;W2W@WdMb]f
3A:JEL;3<64CIP>c:PI^/6^QM37JZZ#PcJ7TIHH&^;69SW360@)4&gfGDeNAZ2]L
[99,@8c)/2;A.6;]NK[<?GQ0@(6+.14V31:fce=UN5a2,QRTY&04.,7(g)[^N+:R
DBbNLfCPI4EP<GRS)F989Bd3#&#ff4DMXY+e1D18BO#f+RO+J\43NAe+&OLUNbSZ
Y<N5Sb>\>Pa4HE\_fWMKBD]La;c:,;,#0,V8U:0JJXS66F:2-R6OPY06LJa+:ADI
6f4?P[Be2UPf@NGO+YIA.W:X=H,f<)gWR&2)DbgU4>A/<[#=85OU9JQa5A#)\;YJ
?-]bH--U5gYVDRVQ/OBMdd0JBIN-PDI&U[_e@]B=f@EUa#\VSb1LL.d]6][X\)@f
T8#L,[gS\C7,JCAX)ZO)97cQ;5^eC-E+\U\W+U>Tc2M:R^a]--2VFXRE<7aZR/PL
S?R\DW[SUU?1O>28\W9=UXYeTSL(eb?,&36<7;0/-]Ad[EKd0=b3-#5?S2,FP0MJ
\V2OK^RHEBA40<,L-2/Aa7g/#E,</7P2A0N<e_3cYQZ>#_f3,&:Wcg9B6<]V7aR,
N7:gc?5WA3cZ90eEKR-2@/KS,@,5X=WZS@1-Z^P:L+DCaBcML0KSN^=T7Z,f,Uc\
C=gMVR[(Y,2aEDLdb7a.MVOA9,aY-f[N-77:BV;B^PGI6]g0V>(3,K9_@86_>6[)
^M5TK6XW[#[8[@(b(/d5[NPS(Fe5cW&]ZeBRB1#9Cg,0@<5EO-M#dceFTO:L#5[P
A.FT)R7^>^28M7A57Rd0&(J#,M4?K3U,G[ab/bMA1GU]Ge6]LFEU(6]Tc]/@B?85
6Fd&P8=;WTYFa+;8fS=I&4<?1O(</PE&0aE@5A3FLC.R.NDBCR?F&R4@4,dUNHdG
K@2R_+SKUDRb?_BJ?UWNQe4]0GBY[Y9=QFG3V[]/gae2+PPd:G>ZE[gGN^PZIXgO
WV&WN;G&D(?=4)\//HfDeJ;81Z9?J[Ng=4Aa]170/d6W=6<55M(,QQ)>JC5,=(cC
ON]b6DIO6bX]U6QF<3Iba,8_LZVA\)?@f-cFCJ_9>?FSD>PH&<N[TDDeLI;HS9-G
bAZ&##7@AOcN?)P6MbNU^NJQB?.:U(L30HVg4=>ZE6#:RUP-8aC=ISX.G83_bTI,
NCe=2NcQe7E@4b&<C3eEd#T^=2R;0IX@XA#IZ9BR3?>;?6LLXI=.@&UC)2EePc=N
J?8^)gGNFWeSe_PEF[6.+MVB\b@g2a0;VDJ/,gY@2X;QQ/GR11](AZGS(Tf_(P^=
A+U:Z6Z(M:J;6bafM7@+_13,]Q3J4G&_EKGF)06g2S6\L.K;\JS:F);4K].DYK=^
g?Q_b_1(@&[MeG/JM6F^R_;7X@@Mc5=K[6eKMATcW3f-CPI]XY)1QcM/8Pd;TV()
09KZ_(MXeRa5?Y^NgJ@N0#6/>M5KdDQV:<\4[1E7>8C;I-=A?^>C[0Q5_2Va(5Xe
DN,>EX9[g=<]gUSO</OXAA7PgKcGW4K,<?GW0gf1=/>K[eaG.IS;RF.?[G98C=R;
D^#[Z2+8GE]?6(5KJH-L]>5ERQ6D\1b8PQWJZ2_&>-76a,OPT:IG2&c1DY;@CBO2
Z>3V2@a:1ff12Y9/Z5dZ:XJPE4=fPd_X)YYN4L[gBI/a-Q]&A]OO/<1HH^E0e77a
&1gTWQ2XPQd)4Q@]V@<KM5BLL8WDPK&8[]QbBKeELMbZ#CH?,J97<5bC2PDGUOg>
,J1^Z.-O0K)^WT@bN;69(&0V-W9MY]C8RR..fVb.7Ae-Z9D;/\9f,FbXAcE>.aJY
\GR5Z,D[PKLT5SACNS)4=P>BbTDf1SeW[;QKg#V[5L>6X((EPN&0UC&@V@cLgJLf
O)7Of>L&5,F##4.&Y=Ma#Ifcf_.=GWNf>(SNL7FJ^)6/a0,gS]^a1Og?MgM9>a#J
J@8[Qd(G&N7V0(X/aFAeNCVRPAGM4(UC[-[V5dKYOJ,N4I(R44R[#S7/Dd\&??,;
1RTaS/3:P;].\CG:4.7:7D<JQL^DZQL(QQ]E\R/Y_bTgK3YGC?Jgf[C5YO9P]BDZ
WS<@+R8WD5F<fU0/,L<0+#P>Y\BW\]DIAX[\.G]Q/?63aH7LZg0X26XI:HXf1\Z9
2>&J+/dE8cg@55?H/_7Af04I<HY@Y0Y#?@BX^ab>d+cEUFc[;9PDc(E:[O9+QQ[e
VV,VZ6N0:6)C@#7;1TFDa][(bWDXMAH:AJZdT9AN5;8(7GW)5J<aRb3H#&I/EI3T
H#F?3G//ZG[ET4;Q^]S2\K.CPJ(VJM09U<Y^ObS9EQ[V7;SWcGO(JRB.,)<I:GE6
W5db#]&1Lg1B&c)@:@BB?V5G5SXZ2BFW^6<WUZZO@_<U,6+H]3SBWV:G?=R,UKeB
(cU\??ABVeM^f:AQ#3<2^aZLLZ/O-FX9WQUIe&BZ(P,:,21I(6Z\1V9YH1[-Y/\6
-f_Dab]fOJ(a&8QU8f1?I]1NEdSGD+M?T:FA6.=,3^9a36:I/?I#d;5?,_>(e6PQ
?T88RU9NXcNaMZf]\QDXI2_@>=#[e^5JZ3@_.&I:CZ1#<8T9/I_^FQ@,19QbaFJ7
f0JCde];2SeDdZd7UILFO[bC:b:Z=gc_D,5>,,D2Lf=^cagGI2+_]H+.HBCOfYW/
?7?&-1CW+cL@\I-e.[0URIMR,)Y71/c.1<\^,++IZ/6]fP6(;P,6DR-@\GAggc8N
b@PVa.f\94LAeY+.GMV:^KW;;-R?<,0X#f;_;OP]+@C9HG-.4gb,K/bQ[dR7F#RB
gMH?D==KbKUNO&a-B]7fYAX4<39e[E=KdC6@QZM7]J^XfFSWMg<J/4I9NE;;>XN/
\O@CL@f5;;Fe7CZF\(RPP)BV\:S[(GUOdEI2RQAI+31/<WC;NLMB2=(CFDF)EeDW
N/,80OZ.G<,9Q4QeX.^P[=Kb9f<,L7HU=0VQ7^-2XU/U//;BHcH2(I]RdJLT[c(G
.JYB#1KZY0MR.c_R7I<<32HUJRJ;Y,ZZ13^7b>@TGNQ[4I0M3a+A0@GMW1L>UHHB
6D_YMCUbE7S6HbDIQU2M->=#bGQ.\B(+L&KeF=ZMgK-8#JN\CQ1@I^8T[e/>9)(B
MD&^_LZR,[I7cL8bJ&AO#+MN9MXXgT/4U5-c],/fG2-R23_UHTZ<d<SOL<I<+HF\
.PeZ9O8CK>@T#TPB@]MZ#E9ef<L.3cT(>gPg\O<;)1/@g6)_69eH(DC934:_RE9f
0bN.QK1aEa)3L+Lf[f,,fUEB5D>=LY1KHXfZAcL.5.C\BUO1@A(\+S&@TJBf&I5[
[WVaDOBJG21>,?[+/0,[&afdgX_g^,.?&e177:bIf<C:-5(DdQ-^Vf++)),f[fL8
KNPDS13IO<H.,IB4aPN_X3C4bW-?Y5M<4;N711L#f#@.LS.9WNb0bS+V<37_9MJa
5E7Hd7HJHLAd8F<-MSK#WXE@FH?W/3gZAYf#7cQ/=;M7G(9PcSG409JBA_6-fcWP
L/4^1\&=5MMAIEQJRgg0P&Yg7@eAT:BM]dI^K#4<V6FaC],Q+#+CUQ7/6>/=IPX8
:X4GW-[-#<a+a0=Q4dgHSTKU<fBFJ=3/Z65@:TT8gR;YE-Z6+VS2f9cHbM_RL;]K
(8NZ_61d12^MU50NZP+X^6.+/<fUQ0LD0SO5a=];:2PJT/ePe1&/R#AdOH;?K9_T
L8J:@B7)68,6<+POQ?=8[M3Q)VI[PDY6>+V<:5Xg&L]_@HDIbLg/f4Q@F\&2LO#;
bYQG]/-RIf>MZeR<bJYD\+431W3FY;E]Nde1[4DSFE9agU@F_L^3.RVPJB.)B^>:
^2b\cSV58ES86JYNL&ggd53ML)]>V-N1Y[97V]XPg6gY=[eHKLS5^\E_=&HV&AW2
SAJ\7U8c>\((6PE4X=N,T.;C_XIK\(3XT/7eGDa^ZWKaD0G\,6GYEK#X#d##^0AI
X2XH7VE^N/L-07L?d_[MR=UD??b@(+MV7MA6,S1/&#&@YI@/@0Ae/YgT?6/A]2@V
HP>87<2Of-[#AX//I4<7FBI&:7W[d5g9MB8Z#QCW.V^:L.;DMHHgXP8B=aJZ[G=[
Y@O<Ng)Q67([4T)A][_S<,a4-f4_gb/e_,?,e0O_ETZ.N-ZebRVFZT7g\?_LF+X(
LQ@fGfE+(Ye07P/00-8GWS+ALf23e5=F^d>BM?;e8@NF@E33.aJ>PBBI.A6b5&UV
T=J>O1/4]7PFMW:)G[S2:X1])604)R^fc>b9Q=PRA1O0WF#4/A#K9;L)=aA02C2(
<=LNe\]R,\CO-JQ>bdB_KNFI.&QO0OM6BF1Y^M[)fd=Yg]PZ3/=5HTWb6D3+.TF9
#?g:4c5><UFa)-0LR=7K#(7>BQQB3R-_&I&ZJ>6O>RNO&=<,+._,#W/]bAYUM]^1
@Y&De_W1<2EgUM)Gb\30:?</fdVX^65N<b;Y7K_bdOMC:6L6ANK]d1]HeZC#/Q^O
HE0f1.<1UO4FKWUA<W7(?+..R4@Pb;ZY5.T1FK(5QeeaMc9MP8\\=<ZW6=]_eVS^
)Y:=:b7W@A4bf.c&((1B32,@/X\-:&b=F428UV_B&2S/I&:53]7P4_>4OU&L8#O4
#eI9VZ<Zf^.WZfVEBCGf\IbMDU5[R_9_//ef+_ISGYW=EgULHU3)HG3=JdY(.XIK
/fg3TU5]NUL23]#,g3?X2U]OE-:JD[\S^<V:<P)&c)0O@a(<4bgZ\^WE6I@aa87X
@&6<c]>764?QQ87d5Q]E\,W05FI(7FBETb;+FPcODbRVMVKeWF9W8UGO].V5eZKM
,@bdG3RFUO5JY;B<82R&,J@0bNR<b+2M.8PAB(NOTC]:DgVIH9EIZZC:DB(WB0bE
HUg[fH\FbDJ8.>NRe7b.YZ#Re6QK59;T7\HL2QE-CD#U@]U4?B7E_VK+Y<47QIJ>
UO,TYPGN6(+9@#C:gR<]Cc[4[QOOG\=S3e]MO\fJLXd@S+.AN2IQW#^,3VOTX7bP
28NdTG;GFBJF&T.T;<,Z>A)SM&9Mcdd=dH0LC)WZ#V-::UTL)#eJ--gg#1&(E+)(
];_;(f^e.]a^[Q+L(W.<aH3-gJ<C&X7D:gVP2f(;A=e1F]dLCK0G7TK\JX7c-9[<
]:@A&@N=&9E#:(P9<17b=OD(Q0^YK@ccF-ET)EJ7)C#E0ZeX?@7>D@7))R]APKe4
-1R0IQ^QOC.Y24C6NFSG1A.))T,\9-O&C]>\G9;<Y^GZS&;O+=MKZ22T_):ebEZK
IdG]a#fM<H_-AR7MbS5EMORZ;CYc/HV)L2VQ)Ha:<DC2W]1Z8)&I/Yd>[C<cTD+>
,&<e?),#C)cg,g41Y5T]C\Z>(bGY2JV)8=Q14Icg@[f,N<J].DH;[JbQ<]8&H4gf
7DfN<&gIZ^?1W=@_)S,N&FC><;JfOD#<fA=8G@E<455V>Y^\cOE_b5KJCPADUC?[
7[1AP=87TbY^4+_\P8\XMI+/2R5B;/c(I+HBCX81#1@1Re5d6F_Rb^KFGP/.JM2f
PM9KG+MVcdW#ST86A0UDM#+/,#YSX^8O[X^;(LT<KA[>]d5UM87U._ZM#=;J-U2>
F<+Cg:XBcJMU[WLY.I;f@.[1b)@W]?D]AC/)E]MK20P\9b9L^g\dMKY.0<@ZcdQa
CEK\H(=M+6\<@G<R7>@:HW+=dG/@TbbX32)N6LQ68]22G_BNXM1&F1F;f=fQY2g9
gQ2CP<@H[4]BMVRP8.a>f->RUV0Q(PZAA^+DFMI&CC3eHbQ1R717&:\dCM;.JI8;
+.gI&@Q2HL(7W:UJ:8)4]_P4O_FaYdUFP^;U:C.L+-F>JA&+NaMR8>=F&7;aS7=6
DLARWGdRVYN82EAV,dE>,X3ZKYF8U=SQ.fdTb2>EMH:cTP;>D_,6M:;1Xf,#BT:@
V)1G;LEEJEDLBa0&>+Qe<:S\]AA#A;-0_X5]<,UYTaTKQ7V/.9#JYK7\]_KdWT&M
Je=YZ[d1c3FCOVUO[6Z0\-5LC&,4>E_GHHMBMB^(L?=5TZG4;4@1Pa@Sg(@R-Bb#
O#J6_C/9aS3AO@ae\]UfTL=-9+K?Q9U4dDU[\.Oa@HB;f1O[7RC^.G@bY_e^,48\
@#U.:-#1G:a/@UHb^A]gfL5P1URCg@0(&@=OaB.&4eTW&WJ:6ZDdEA5_G;/CM)H>
?VUQcDfE=aEAOHB7dT.[B5G_B^gL?dF8H-a1^<:TM+e(BE#GWZA3UXU0D[-SRZgG
D7?O>@G>]GDWNS-Z_^K.\BV\8H.d0Q>Y51:;f6A2=NEacOB:Y_:_HGLRcDF:EXXH
P7(cJ\&^ga5N5JF2TXM=Xd\_MAJ@@J^efg_HX&?B]7PfN/,&=W.1fQ,TJde)(^W4
7W).HL3NY0Nd5CM@JQaT&A5dL<;R8Je\A/<^Z]1eA5\6E@RV;<(8Ca6.@7-^bY]d
-aS:cWLW82ZE47T3\C]7,\_K7g8g&FRg4U]A6V3SRR-Ie92XA+b>Y8GMPQ:K+C@[
X9PM26M?+5WC#Z<5C.:O;<DRB3S23L4eQT<N;KD&3<X7F17FITVNODB\/g:L9\:6
]fJ^=HZC9(aZ<bV@2MJXDII_b7&95&TNT+=6)=?;\4BJ40,^/L2bHcYO>-+eB;3X
?N[E\4SNRHV6<J+OHR_P](Jb(c&DQJ5(a5_BFAT5Z4=\7d?KQ^1:Q20LbC[B,V0d
V#f<9DRWERZ-QK&@R>aC>O&QQ=&Q=B50R+4FLO+JLXAN:=F.B5[UW7;;&XZ->R#S
#,#PK<Q+Ma>Ncg:S44XNU7#Q/K^,6^]T)5&aK.VgHe5a)NCCb]5@L=1cUR](>YFP
Nb^O7_ZIMQQ>9?[T]>ace--b/\+BMA1:WI.7L1cAf&R+C.:cJ/)8f?_Jg8g9c\DK
428+EaW>QbOS3L0<U?74JZXRJ3U_,8^3LXXg3S-5OXZ7AI5f;UL.A37^HD20AR6I
c2&5=(^97[;8S4\U.-)DHa?-GMS:JFU-A&H0HF.bW<G?dE[f]Z-+M^_C1DLeOJ>W
T)0..cLEYIC,8S+&EPSXQbJDMbMH>Bc4FA5dg0#@P\Zg\<7H5XJcG,ac/I21&]d.
4B8LaMPNPfV3AM):e>Pb6:,VQ@EWd]8.WM2bT7+2GDLe2aY#@Od^^L8_#YOU;RPH
R_SK&Fb=3=,c-J217)YD:+\QD/Q-XVDI]CE,(B;c+I^AdYRWE/CF,+J=T\Q:_6TL
G?Q+VEa\I/7(?8#88ZFg;+9-X&3(e60JV0?cW:1N>+\T\Q7cNSA\1PN3TS9VBB]b
N.SFF:cBc\/JP?L)L#-(PLWP8NS+.XOI?bP0eQ\G:3.]f=;,8MA;?XX&Q=4D)KNG
P#U.5H68?Hb-AbJO(c3]c)VX4^WP+a#PPVAb/[f:Q275\O(V3;aAQP>D;Zd<4ULX
^?/6c^1P.O)3#^YMAAXB^TC8O3GO>,M.GcY(=D7=:J4VYc,F5dIKI+;ZU2M&4V#:
;0ZN5>6<8<Y#0D1NM9YZPaO@C:LK^gM[#IM4]/aXWY55L^.LeF<K83KW-#^_OfD<
]Lf_?AeK7E[\bM\egeMLgKJ0=K&(a)U.^#^gT&/0?/3#eHdP[AX_M^P,M=@?75b5
>P_#(Y:a((^a1QaSUHW>DSF3,CN[^J8W86^9W-<H#W/<<-T^2cR3\_KS_1OPI@+C
TUYAdU8XM/VS7\9V[74<b_>+a_;/\M1S_+A3g-H@J)##_<fa->&UD>^OH&Nb;W<f
-Ga3<gKAZLN//E3=HF#O0O+YCf.V=Z0)):J(FN)SJ7=A\(E6<Gb](<E5GP9FB):1
=FX/Y6:_115IP07-,I0J3)&1<_;J#4;NGFC>8/+e#8U12H]R+_b-U.E7I/]P)CP@
#g=2<_#V9#cOAF>[3NS1G\J1=@Yg-\F6?ObY&AAESf\2G]99VO)XZd)V61eBUV+R
QaT.U5[Vb\M_MIfH4MFeXOcH531S]4JA>#DKb5]B]CbdZEGEQ#WcP0Gd06K[eCf+
Y6KfKAH0FYO#V<a(9Od?EH;VWB2TM/&0<KJPdT@URGGAe;c1),K:2fE6e5\XNLQN
W@GBZ2Y<\OO/g10_af16V[&Ga8IYL;Z7VdM7EMbIDLHFHdB3Z,0^O?P&DF,U;[-T
FNZI7a<7+<9eaNgFG9^[-03MWD^KFU(^&ILS#:&06H_a]Ie&_LOS+(53<,H&gLW(
UY>Q?NPXI3cSPV2[/_6U+92be40],5T9O.#^29R<dJCb^WX><1HUb[M/;8YAZ]22
SfLV3f\0W&H6QR:d,7:@A9.\C/QCZ&g-NW\daBfPM^,V^Sb>5aO33_&D:,J[)g(.
9c5ZU;8Y>>/LI+KHC\F;I-fE2BA3-(_:Y?d1Ube#?MI7-D]1S=@b;DM2GgcN1TWE
>U9LV4Q__e:X9#I5YD)X\?DAfC&&=4(IEL=<XaJ5=Qb1Q5MBSKX]V[-X7Bd5J(+\
=;^G?TVMSR)Q1Db-LQO#PG2GC8QO9dYB>3GTCJOEfg8DUVYgKMRb[f<]L1W]8GYP
VdE6]3F[SFGH_E6.=0g<Q@bOf[:Y(YcW=9MGV8bPK#SEK;cZ:P+@-FL_d7B.]D+Y
=WbE[-^IN82+^4d6,8QdBZF<<WfH6@^#M,V8:(L5P0AH)T.:g+59>+8K4+WdP@./
Qa@+Zacff>:Q]5D&[?:3-_<c?1>5Y\5QKcHDLOP5VX+6O#LXAJ<>I]aV\0:RQWR5
M,OJ.Lb?eZOU^L)NK3RNJC?J<0/3R5H1W=@0IgAR6\P8O7H/<e.[bgTIEbW=3-PM
:Af1,J;&Qdc#=)+bI8G0QJMT^cfZF8R:[TPID=AP0;f7,-Z=8d^X?OQS73/DT7)K
fBBK[X<:aGJ_J\T2YOO70CH8aVOI\_[WB=31Y1.gG\NI40^G4B4P4E8\7f=g,d0e
@;)_f64HWNc>:PJM(;KX8bM(S8=PG+-3AAR+CabB5@W#BZ6\+d7<c?e/6V=9Yb/S
J5NW,Yb+L]CXZ>=OD0<0AE9NFEU&(c]_UQ:d2(\bX6Nb9+K]VGUC0Bd\Y5Q@F3\\
7,PI.1;?<,3U[)7:]ATO@J-[1-\^]T+B]H-=F311+eR?\g8(3?+BG9bW70/S=5Ob
D=+:-[4R]HTNYF/:ZE/+(LM[_?bV]C]7+LTV+9=C@\A2abg#0+67E3QXfN6c6EFS
F<Tg5H,IC=SCS4Yeb#H33_@ZVN[+O5bg4Q(Y1L_W[aY\^3-.]F0OQ,>..R(H29JC
X^MR=c1P6=0R2ZZ/2?Y(>D><\d-&TQRE32ZDgH=;AB=F1H2[/<P?2\g+P^cVHaaW
C]CR&OTadddbJ]?9D<S2[S7<L#59E)N)/+0/MNfcZS=a0<=+P_0TfPR=@;?.28Yb
VWa2L-0H7dbIEH-4H^D?SY+=(@;9)@Ic\If;=,cEOLKHd5^:)ATF.6VM<,M,Pe[R
c8>;cE2OVgU0M1[Od5E]S2YS#H_CT@AJL#549NG,RS?f5+\P?1/4P\9[Q8f=U-^A
BVa(H]P?1O=3d;S/W3M26#8aLCf2adRDFKGFCV1NWBdgK2/WUJG4=:7W;;L[X)g^
GB<abf<Z;,Me2]g(PLL^J3>?H.ZX<OKM+PO.4=3<?Hf[c/Sf9.,)-AQA8O@bIQBP
>2g.OcFD9Z30H.6F?69DPF_6a8AA;>NQDH<I[7V+2N0&U[JE+<,B;_]S5AW9:+gP
XJVH,RJD,X)I-Y;(ZZT81:@TW8c),#GO_Q-J_QM;NUJZ4/bf:4:8AeN)aH0Z42D/
Z>:#7K#X:3.2bO@4>S5C5\]f@dR&F@fPdb:/7QO;DF[/1e=IF:5P\#Z0Y\8>G.bC
=I-@+0)M1/RCD9/0BGfPaNaGJ#ARcMeMAIH>\PSZ(@/WYNdH3/#4V/21=/;UV7O.
#a@WFcG1^EG<)d5C8)CYLfK+,\Z[K\?(<[FPTdX/^6ASe?\Z<KJRb?Ge064V00B5
NG](M=c(063(1JJf+AK(DLY-X1=F<+HWG+,gK/(R/OKJ^R@7HaYTL7]&UL=)MKU(
2f)+Yg2<Y[VfJ9O?)(Va/H(X_ILaK\&/YB@0@.\USIHCR\RS^TF<^+=TO03eY)]>
,,C?4<-5EVb8/F-g2DTQ=R#PYUFa>b^&_e[<cb_QCV25W?780C\NZ@aP6=-d5dIV
.-O<X^39TbO[FT8@1F6O=IX9gU<37d9N,B\UXA_J.(<Hga^)7;OF+9Eb6cLG-_E/
SD,.;5N2g@4A8+U8cUW:?L-A2)-WN:YLST60e/+^6+e6T?:+:2P)/AeUa@Q0Q,=X
\9GSW#RY7V[DATe=N6^L1Za>338E:e#2PY.5YQRI438f5:fHEW]CX2=36Df2\bJF
1cgB@5BRF=3<F:d6TcG@WR8VT2J=S_26J.,?+,-?cM;aX.<Y<7F.1KP=6gEd:d;<
8+TcBKYIU[:gTX+0/<@gEaJLN;3)&G#E_B.Q)PH=F4@X/SQH.OLIKH[7+]D7dIGR
4TKJY-ZW;YVK[&&F/[cb+PWA;O4A(=[DMTeUD/;D#[T18?ARR=N05[_N1.d?2+61
57+?acb(f)d=1>R#<,+E98(X06CNa504UfUD&U3Q47U;b.9KQ>:;.KQ8gc2^@UU.
>NDfZBAOeO664IB&^<(77If7cSGHDCGb<QN:9&>d/F1?V?I7Y\H^^>?,]B;I<#+H
IdaAR2f#]A7R,(@aF05D&P\)S19#,0G]&#W]^b&5YN.C<QI7./-_=/._1/R=aXU]
>PeFBK7RfQ;d[T/2CBG83-H(U,)?\,(#EX+3F,_0SaFAg8),]FA:=eOO5ZVFZ1OM
6gRAOV^X=VYe,Q7g/b6<c]N(E:6=1^AR\cM&@S;gP=88Cf<1&;OU4A<]_f9A\,&]
V>EFN]SRCDB@F>bf\33_(C32I)7QRUe/GP7INPZ/00\Z>>77A)g3=S2V&OP#/2YP
dUg9EP55I5B[(Z1eQc^,gZebbd@_(cVXKA0Q^]#Scb@KKAQ26J:?[P,C82(XPCU;
PLc68fO<LLY5^JM+;fA0I\C(K=[f(CHIDIJ61TQ=/Q^,[&Zgf.233_PDM1M#=2fL
1@](:IFB&IdMSQ=YCX5T/fS>&Nf>Y5E:WKB<6/aY/M_4XK\9L8?RSQ1.::ReJ0&I
)b<D3Ae?ARa+f,#_X/Wf;(.V:g?f>Pg:TAGgI24@QIP]UQW]D55PB-Fc_bb74Q^c
)\1JDe<^HWD>Nd?#)g>TMED<c/QcDUA&ZdH+.]>^#Q+)9ROgJHVF&90M5I+X9+.)
INY+:N3EPMd]C.B\QXJ511(=ZF4CTOd9f_\MM)Ja+X098f::17MC,d]Q0CM2@Xd6
6@0H<(42<1(=7;D:AGG.PK=R9^B-,#B4YFMT]d:_O(\)?8?a8UZQWa<H_@YR17.T
;Za:f]GK+PAF6:W;I\\^GHZPW[+@eY-C71WK0ZT?YBH[c=bFbd]&GC_U5./=6PX7
c&16/?0;UP-0X+;(HcV4::\E8)3J\K1g&D0AQg]#-?\[O34N=.[SH&Yc;;XPD]g0
KbC1CcL\_e7ODV+4ZFLX?(dNbZ=U\O3@cUXf+O,dGGfI^5d(\THS;Pg5>=02T;1<
4GGUT]T&FQ<(_gC2.XSZbbM@)VgTJdE3T2K._1OJO3DGVfJEBL=AVeD\C)]A3ZO7
-J0>Yg+X8Y/N,)SggZ(QO3=Y<e6BN^G\@W\gOT[N:D?SLL>?>dOU?<XKG3-K;0<7
-6E=gZLT(RLLA5QV=F-7QK&L4:=6\dH)0<+#&aF2W&/2SF;[We6aA__0=XC(ceJA
9RO@dfJR3WR\?+D-IAd6G#=D,.&[)W6HG)RP3W(=MWO.W\=-&#X6HS-=/@V0?A6:
Ae>7EPW>UXG,.:ga?f,QK8>SWF4K-FEZ=cI&3@7XFW8PM?&9L5Q@I=V,TSE>M.6O
-eb-U<SF/ELK<CGd/QU?@\SKLP8D=,UUbDV^Q@D@_C/&(]J]<3[IgGg7&CHXUU3(
&L3FX_bBIV42PRcIf62b6Y#1cY/<NTNOe@#KN@8KX-0S])N2=C.;4e2TZ?L)T7JR
QV@aSgaM,SZ=YEU94ABXBQ;=B6>VP5H?4gFY@#4L=^fQKJXbXQ/bI5?,Y-G(KZ4]
5@O:YBW0?)=Y-S21M[&4K#0,fJN+@]^NC.ROeVG-9Pc)LPCP(EL0Z>BQ-:ILP8MA
XBCQA,^+L5_+U1:/CKdJc3Ff#d;=BUM2U(S]bKA]/SQ5F[adIIF+?=\gS&X74eaC
^;/d[H=_5GUAB4ALS,Cc5c^2P-;/G8CE?RRR;dOQS4QS^<M\ZTQ8XJIRO1a89bdB
0:,^\N^K0,/P4^84#\)LQ:D/7+R,U/OVV<2.-E&BaU_WN<Rf<_(ZPMB8\\Q:8[&P
0)5F>\MD],3SSYL(._a8b)S.+TEHF4,eA=RZT:-aMM9DTSef\g10=\PVG1;a[D>9
ZZg#>Y/(IMON:S3Q#OZZ&,CUO#Ue&>\5/@=-26Cb^#Z(dT.P@S+]E\.HEHB^C#0_
d7&Y;W1(L@GQ;M](S@e??FT6d861JGL:UA)3W6[OIH/)@cS8DLdMEV,4(aR>c=^;
U?XAeQQD,VRFe\191a#UV7YA6\YV;06+IN6/Md2c;..@T:OE&-B;5:&bW3Q^<WJG
I<B0baQfWBg2H+;;[X>SHBd>I.]V)6dO6_YIJA/#NX^/<LA6BNVLA?M93QB9.34&
&RBeM#W]GKMW1ZP7MI#Z_::2F9]]H2f:97>-@/>K/dX&EH>.>30-2O5<2AaQeDR4
,C3e2daPZ5#@(N64LKMW;Z&YRaA#>^Cd58FC([M-QFD\3L9(;/WZM7F44aEQP)=6
P+>f/O?:)4F+QZJK6M[)[<T?;Ta390FSa]+C(e3C[\GUPMLU\EY0L?[AOU+=,+EL
\RA,M2+?f]K[74[H+JLfY[(cF7Uf:M(Y&@0-g.X>LGL&cgX_,TV]?N/7N3f1\>7K
PXE[fP_=T=0W7(>O;8Gb/IGS186-P._be+f,c9[6)K,+#EDX2C8G0,=).VZ=384e
4KeIF/=CPcF^<B4X&Ka=LA7d^X^MIRQ8RdQJbb4+E#ZR2M&VF&dfCA0+6=)gI]d>
9Q<B-5NdY+#K7X<Y6#)@:Fc0-eA_.X=9Z_:W+BN^7D_=e-?:RK-LCJC:Q&?/O06K
-@\H-PO1:Z7XI8FL:<-6DA+a?WO=R>1)#L=#&.E](T7.VCP_f<Wg>S8YBc0R97/+
,)cJLJVN[01[,M0#cN(FgW_@G6AS[[ZSf(;REE=X)Z2T<RM&JCJ(3gEa]S1&6[I.
4f<?Jb3,L5BO9+#\^ROC&bU>;[2#Q,M7(X65BCTTQW+d/(gD(CT^9,33=KcQUV&D
C^2RCECT59W:?#D5,<HXDU+#)+9G4U\C,gg2\IQ]P3G@6d1[?YDb)Z7_,4+\;2I-
YN(aP@7DV0\:+FRV@GKUD.+K37Q,>a^C\;?deWAX(7F0GK3KRD7_43WeNS4:U_71
g@NFN-O@]M^\4?1^H9XXRf0-<DVgZ#?[6F60VbS@)5M,5[PBVI[=C?])[GR&fR6,
<S2D(?K;OS]KedR9FU8fa:P,FP9#JYWaIbJg9Af].)F5&d:6-^3VZJc-fXJ4:GH0
Jg@@X9c10Ag5#eATYKB]dGU#()P5T\<c&R?M@f?XASg[gRRGYV6a9P:.O:L+d_VR
WPAHd+P48e?:Ua>\,FNf04J[YEP:W=FD,a(NGK(XGf[dWU,WI0XH0V<FDJL1\=)W
LgdNAeLd(6AY0IbO(#AB[F<T(ZMN[R4ea]BJ8f/BAY0-2MQICUb)T#?_R\,c)558
F2JKC,-CDT1XZVYD1K2H=S.TK,cP/#CM5LV=ZeQ;GL/VNZ8K[]b4PYVI/e@H2)RN
9fb8e,^BG>+.VF(NMXg]ASaJ2&E@0TEKW6TDfXdT[C]GH9/KYTIP/3D@T@\>&fc^
W=^W\#DeXe&+NQC#NG#/KOON&_8\HBG()SJ4G<V/NEH+BU-+(^ddV_(4^678W3^\
S^_V?FBXM-2.1[O1G>-N0aTF4DB+)&72DL(KaV3eJ<E,R34?FNJd)eDF?_HJ9Y&]
7W)[e0MXDE&XEC@KO.a7@b-42]Mf2:R7c[8B,.7N6CY\-JLD_S/4?3NQT[M>W2-B
?,GEO&:P)ba2>_DE\[B,=E#8V.g>5-9L.eWUKP=O68-,<G:)16<#U+eNLV:L8#G/
_0NQ;\>QGZ.&-W2?YOV_3VE.3Q)/(TQgW<b2@F,B^5=>&L<5R4:HRJ_+HD7^ARe3
,_KL.#/XUFH]J&DAQ6D?,T.b\N@CS,L47:,-a\dQ1Z_>O,XZV]VJJ@MO>6+c88e6
fMWadHX3g8#+,XE9<>PD7HL@Ib:K)XN3&=)LS(4c:^KTZ(f/67OQ=27;]T.7#KM9
PZC]#=V7A/P\W7KQ>:J2TW#=?R.TJF_=P;:Og:4=;e+B<^VUa0I5>U@FM^ZI+bYa
bXcK_b)fOe@6c;J_2Zc:a_\ec=;T)G250P3g)U@KFUH?aFaTK-JW^A(KTJcWB,,K
H;EJJT2(g0]MXS/]A]J/3F=?Gb>#Xa[CM_P5,gO7:Q2;<C@eaI0aY@/@^KTPRFSA
bW]P?V:G&c>.eMK9(&3E&^W<aH<BG7G5f0+>?N&#aQ,SPfT;481OeB>:OCNR0=3S
+Q;9>[FYe=YQ>X_9]:VVVFH33fW,cMKA)N71c87Q28I1R=7L6QM89/7+:+dNU/#E
17;9EKcc=aNY8=TIBb1/K+2AU=3aFRGC>2\MM2_P>#.C]fQ+W9^.O(SO3-DeT^c;
J,)dAa)e,aK789caO?cG)1?f=_dg2=(K4EM^Pfc(@(X]N=[+E)QVFN?MB/Z>UQGZ
X3)cC;UT/R;](SRO<CI@CX@,b(Tb9Q/Z/4U4WTH+C<Nf;^\BB=LZ^IcMY)1\?77Y
DaMG4\AN<G39)V:]f:6OYYKOdNdc)=T-Cg(C+8-8O68)cc2LE&4ZH1_2TLUT3T8I
[5bQBN>8f2XY<ca/_E8TD#a1V=a64?UIX8Uf17BS0<KU>X4eQ,I7OXLb>Mf9PcFD
TU(>AH&[J.?R#gO@&ZSC_g+>L<OJY.UJ>a/6QeVG_CB\WJ4>4BJ+3EO(SYC_OF&Y
9D5/;<f;eT7Y^VD9WWg[_6+HK<F+^aP(Q=7(E(01?KGYFK2dXZYI7V-KW)P.Af,Y
;UEAWbE?^R]V?BUDg3)CR08E>R\735\1YaeOE_gEMf0ZZ-ID8ZR7Q/I;&aFfK,+8
c(d/P=eE^ZINOJA#M.O#9?7eT,.XgF5\#/5e@]DdVag\=V@YCF:XV#ZIV+]P^CR+
>H?Q3QP.7>S@1XR?VRa4>R9&<&X]2LPT7:H\<Q5/S[J5=^=7J@<Y52R38F>LX/bC
@QGQKQO8()UG-.[YQFMcL<_/46aX(^OdQC82>e#S5YXa=HJ@-9KEd(J=#OL@B&EE
aZ8\0SS0a0[g6^DTEUQW<@3Q-TdX?=c1f_(W?OKZ:V5ICP_CCX>DOIZ8.H4@\D.b
7JebYR1Z?6I&I+1QT3V@PCdB#N=VS]6)2/@^=E4@5GN-@@[NF8^<+/3bW-KcDcPM
U\&5OK]c1&EaBZJYZ]L.+b5d0g(-X.4JY\G6+f>^V9VU7P:H<(EFf](T<6F8TXS0
3ec/\gT_,OPUJ2FdQ)/]BgX<N)?JeV?4;d^S+_<6]Qb.aPCV1:=KY+3U9N@Je,=e
J.&+<KT.8?R80^AC9:bKEd-2;cY9PNGd,7YOX]6SZ4g<aM.KQ1^BS6@#1@_?RW5B
[-+EY-23C);,>(9Z8KERBfd>f7SZ[LP5-8\GK=#N94)LNKY6M7NOeZTe@OV2]eVR
(2,H6]06]?N<00FdKT<0Ccc9/=8T_5?5W-YR._U3dYe@e=>b6Ub<15PCG[-.:I?O
2a.26S1]SGeK1@FC\:@B[BD9fT(?)Xa;D?[c,+.+Z[EPN6W\=_8He4<&])aF3&/U
9(T=<89D+7KP#UaQSJ>(BWeOHFVIRN63FE2Ae@3FK.?RUU?\:Z?&P^E7]dPODD_^
X)^?Ug,GJe>3W\ML]eC+bZcfA:)0BB:W8&S&&<HVX^\GSG)=H6OLcJLZ_>,2(]9P
:K6VH=3H#DU0H6#/fbO:P2,g4>1B(@-EJH9^=Y,]\fX03+<6@gbK5>>&GZU[FgcH
JQRJHSM[8-LYGGb/cEeJQHMZ11;0a]d/N3T?7b,FT\_6)/XRaD#8\.V4ECPTVN;-
>F0)>^HW]/@D5VH-Q(Y=:@>&/_,/_XGA?1FVPH^;?HMc[6UP>Nb^MG1:F+LWc-\X
XD\[P35GT6S27BB@N3;P+VDX&\T_9?a\=.JKO&<fdLB3BT_7abK>Ice)e]T>&O-:
9C58&P;,[Q+(N(FST+E2VM;_1&P.6(XL89Yd_=d9P=C9B)F=-d+8C\Z?->F;:DHR
[F?#_)D/4f1L+>DR1:_1.1,PK+^[ZDId]WTT_;8bO2JI[6U.g90F[</EN465ZOF4
05P,@Ag.(\)6fVCQ:Xgg/Z\Ka7AQFV^^013cHB3(S=W)?^4B4faS1NQG;74a0V@;
//09?#KI>b3/H;TR3Y5FV,dYEY4>G.7&A\:?WTNARPU@>,Ad&L8,^HM;[<@VP#9#
N9Kg&D9#Wc),E+GN=>7EP7L>X79#8FP-5KX1QZP:N>gA>FL#98X9<]2JM/0S)6/_
)S&).=bfM-S/O[Jf>#/0Hb(:UPWUSaRV-:Rad;/cB>/fV<e:,VC?HR\g/Fe[6^J5
##bSf5AQ\\1#9b_HO@N/:SAX>]10?;^^8)+(F7P]-;BF@NU0[X[MBH5UD\G?:^C.
,c#OWbC91V]RV@JUN,<NCKFN)0<:?E@B3(1PCB_ceVebQW@:,1cg<Ee88<I.JaUV
D3)P8f@3_M;K+D;NgF0-DLb\;4V)E]YXE\<f<SS8XPA1TT#0<#02BUJJ.OB8gNL-
CZX)O2R=gSELf</@]VVR)JR5MG6,D<C@A,S6:0BRg8Qf8+\FIQZOb/)PLd1WA<QK
.#RR.V_R2CYGUFcM39UEgL8>F50(M3AV:SKLHIa:G8N25_<#eG,;Pb\<gKgP0(@8
a_5VCVL8bY,:([7RL>XbLTY]YecS[-dSWVc6cC;Xcg\7\WKT(HZ0T8V&417?:Z]5
^D9??(MDI3&G&]?GQ6-P&fD[cPAU3N,^@Q3QNYDcf,S]S]7G^S_CRYIJEUVa4Ud9
PePJ^)Q@eaXa:G-(:+Y1C\PO0B-P39W=J[-_Va\?K>)Xd\cEg[G?N8S.+0<NFX??
:\/ZYdA3=;3X>#7:355]e)\#V5df3Cd:X-c2_EZfb4Y.=2;^@_cFD6][F;XD(H09
QS+17d,_>BQC@]&>7ec8#L,V1W4ETFd0U[(B7#X?6L;_OH@)(T1T;0LL,:A-:=/,
Q0,]BPSC^K[&.9T2#BT;PgD>1J5L@C^WPQ-BW=JF](FDY]@a5U\e-_+<C9ZBg][5
X/<,?+aMd-.)YK+2P_Z_8ZG][NBLg,:M_#^WZ&VdX&TRdLa[+(7)d8Z=3D==gcWU
BA)3HX2(aSSS1FVC4\GI#(:PYU,@6NXcJ(+B?NUOfG3=<VX/-Ig#6N]X:^V?WYT,
KB4Iba5>M.a.8))G=+7gR1;FH9FY&aUb@BXG<C1fIH<XH/0g6WO)<fJL=d]?b8B/
9TaZ/e>(+[::4KJ26])&6R1cgWQAUZ3[I9\f82W]AbA.\)8<R+.1;KNRQ9<E.6.E
\?18MFJ_0&5;E6R3):W?+a^PTc7fV;_3e=EVg-bBD&(J1B9SfRE@30gXA(Og?>(>
VXZ?0g>6P\S[@TO9<3.E=67?I1)C_V=bORF>RJ2RA@OQFU0;aXd-71QT\13cRPV/
KV5a9^b<.AKA,:./:L6XO9&_eJ72Y6J@=_E7K=BDL-GGNgIF&Z@F5-gDA)cJV;U9
TB_L2N8/&T:gI^9c;T2D/;0Ie:WBJR4\ATZ/c.OKXW[<6YCD#4U:a=cNF8Qc&RY/
D3;<_3KA/ObDCY,-a-<(](P\Hg;G]0<b+[f@S;FX1-QKg[=?1>baf>O(_dMYQ.DC
Z1UDH45JNOQ>1.W<)>^9,9S/-TW[WT=[9AWafCSJdD+@RH6+,KPPI6XEa;e(P9-3
aVS?FZ[_F9bg>(V9NaYGe8\+:Y[4EHODD(;>^caTQP7;N=E0?4XYRI9]^#/.\TS;
;ST3D8F/KMK]5]^Z/Z4-K-GV]F_[[X[e\YaZ[53<\Hg\2)W61H;9]S;F)X^D)+F#
JXAIJ7O?@G@D:@L[C29+RQ4GUM:8#T<eb)1DV6G&34X2cMD,(?9TUMMZ-+8_Xf;X
ZAEbCBcb,C8,TVPYM\6UQ+>FSZ/6&B;?;@TJH#G3#&\D(]_A8=)]-\XW>V6X3C]S
701:0&PT:4A+-/e9FbK^B.e=E]587GeZFAL<(K9KLN&Vb#3c6+@3:_OV=?[:\Y#6
ST28TE]W&fIN#/()SK^OHTHbA[T?@?EJ4\6dW_A:F?7QW1&-N/_ZgUKO/\7gRQHS
>HF3eGH\:^@99&9,HIFOQde69(3N7?6/+0#H#WKD7I,0cEeUgF;]0.EfL/(XT?cc
[<eDL(YFa9a4D:9_>I-5G4UB;;JSD1\9?F])M-YOV3]EdCI3MaQ6/=.g]CP>=JY2
S?4#H&J<(,UY[VgI5.>b8gJ6A6&0&]C_3:)HgD72]?1)/I:NS-GdOb]-M2WVAUXe
dM^49TYI3F]Rb1DAS:3KL_F4L+2f;BE1g=D7#KfSH6,8=7//8+C+Z.>/G43E>f\d
JFUI-<0NGd2A<MA>N_g]]/C0EAa>HfB>;XFBK_J5N.8:EH35<F_aLT&]EYR;T4G>
FDH:2;Ub\I2CR;@[5/;5B2H61F.X0L:_H7M.YWEggaeOBb1CG9[T@0K+5?a@f>A0
XBB,8d#Ed):R_6S+_DT?4ZMc7@P-21&.>#-WIA(B2_H\73fTN&7bARFd:[M9(N\6
5=#?T8KS@[,_/eIN)Z:1(+-.I\UXYdB:@BbU&8W]ZV_EdRG6,&F:b0eS0L60;SO4
(K#/d(;8CGNBb.a?E@ZI7U.-D(#W(=LZ(7IGZMcNJ9HdR9Y,/V-1)^;YK?0(6^#(
fO_<cQdf/_V?NI:>GZ_Yb^0T#A##Y9)A2B3KfKb=03-E##;IXACE_^CFaFIQE&-P
a8gX>gg>XGf=,PQ7DCK]Y-].8XX:50M+=226&RBY<#9d.^OTIR>S6&7^IOc_]\1K
_L.;(#g&9VUC&F8ZYe(BB2aYPPB#PfYNL@DQIOeeHW_@#V?b8O()J#E9+.#+OI_b
Q6[X]KDS5M_d?@X[Va&L07@^QU9b,)./AS1]F9[+[KO=Z3daZY5ZaZZ_KE4T+^Ag
E#V.]9_:+[O#gE#N?[U/d(D#SYINLMV+J1a-S@cg,KO4d>;INU,SIH?Z)g?^51TO
)Ra)[3TUCUPRBBX=<(-QW7UWN?\4LO)M:D0dZGTEZS;1a<dL;>,<Q[RG^#H?HH#S
f4;EgDB1ZBc_1N1?XcX0YE>J[7/M15:3&J.Bb=^4LL=][7b(-S11<@]<f#)Q+WTL
[LCgL4022O(V(6eEa_MOPbQ7MfOK6&3>#7b8KD;W,B6Id=-)1FK]IRRb;A^O#?Se
UKeD_]ba_WA5Ia&LTU+d\e9HT#(-4Q7E,\CJQaIRfNBA_+R80S)YGVAZ]V<M#_KO
U:[e[K?BKX]S:ZD6[OZU@YTFJ&0)U/6H0Jg3gS?A(LfF:JY\,I62&]L&IFf7RR7[
LY51)7KW8:>GYQe4S,N]1E+bANUV[(&Y#e35(90K7^R<C;2FXGX</dY1a^cJ?KSH
^KgNMMT]U^c.CO0+X4[C.#18-0=M,5SZS?KE/V/(GQ:P,>e;P(P92>23X]0M(^JA
P>I2Rf8W2-g?OJ370,]#AaXR5H]Ng[PW.IPN140[M<W\=00bg-L2EH4_e(02DUW>
+NYe[FFdb-4K<L&^9HT@2JC)2&DZ\cR97==6P,LEC=cJTT>Da:[H82E9LTA\;Y/F
=5TAXf?CS<dRK5J7G,X8[JU7>+\NGbY4^:9:BQM?G7GgCH7R[-ZYb)^UYVRORO72
KEOQW0B<aaJ0SeafG\3>(,=@9TKA&;fg;4N.d71+@cW[DK,:T3fPaJ<S?2S2D^1L
W4M\RM(Z_bGHJ3@#^IN7-(,:b7G&4g&8><?1E;S2]QG>3QdY3[+eaZFF@+5@KU+/
-)[;@W:d#+=G@+[\KA77U/f9_<+C175(5f=7&W^X]cW8,N8;833-<+>;T=6_HN^(
&,@^MN&&T5)DN5NE[&/F>+Q8D+G0?;CX&.99ZVH9BJCM>9-,0_TN5JEd73a:eC?D
K_P)LBL#&E=FIbf[)I9^FJWTJ1XEMXM;[FCI];-M8>PNNCf9SDNQdEa&,RW=JNKJ
X#X>T20_fGM[6<:WbK]B:EeAb4c_N#acWC:4+<F#=)OZc&V0HeEK95:>?B[I5Wg]
-(6J6a@f([-72PeF1bBF,NQIacYW1UM=5[.RTQ;M?]8OX(gI\/>B42+EVbRO)L+C
P]3c&\E=06ScdS:Z[CM<P\Kb0H/_FI:c@gLUf(b/cQUX&_=d3_e&50HV4OMV--WR
ZdG)J;dU;^c<JVN2bA1[Ic,EF^EY<dPSD61gGL(_6KeF_ARA4#5OQ_[F&]c0>16F
7K0]O:)902K0LL8KZYc8ZJ=fLg;P.-RVGUcEZQKU()eV7XV7H-:RDQg0#3EI[WRX
Xe/-2ZgRCT,?#DeQdd4]CgQD(>[L5KY+aO)Z_g+IgYYA88QESH=]/b]^LR=R1dD_
W.[@:2;K4RD.f_QH_RB\CPd8AI9g4[CN@BB#Ue+D0KXaaL_&gSB9I:IPZQ51)ZU>
7QgD.Ed<(REdD5H[da2]212gBFWYc,Y^4V8QJQ?D9P\1L3@6^<]DR/V;LfQ+@\US
^>#9g.Hg:[LYH?AOSPRH9]&62JDTMc=Cc6,H#GBgYZ/+2W[<.\f,Q[bZ#:<A61EF
gP3+1]EZKKe8c(WbAYR;Z146g1(1[Me\&NeCPDQ(@M_-a8X75,=J,IAc3E1]7Zc]
[^>a[;#?9&JeIX2KDIg5=Qe=ZXaA<Zag@V4Z[M9::RgAF\^K+1U>F]C9VT-NW:Q4
SY[J/^#^c@ag7[I5_1TfT2-bF&f4^4d2=HPe68aV&Oa[&@LW4MMN=bJY0g-6\#NO
gI>JaEH#PCQ[Fc]IQF+f2?#AgWYE;WM-8H[A[d1>P;4]AZ#g(f8@,^Eg_ZZ6V9S?
WU,O4I#F346?+WO6[<4O0Q]()8=0c[#.bFSb3228>I)?W@RZd)1L^NRY5?;2M4(W
B_1@+Q(Y=34VB:,E/EWRgg+D:+\S#20;7M\S(MNP;7OX^ZgYgAG-HFJM@,==#Y3H
W)YLe;^OgA_DQO:Tf36H:VCF,&ZcJ5.I?-X0)ZV[gEfO4NYD?/:M_3F7G@IO/Cb9
39c]V/0J]&Y<G7(9Y,I3O1O1R:A)Z5AGdeE).gRMX4P<YYP7b,X>dDA#F</?B>>E
3(7dLeb^GbL1PM+f89:9L\A#M/LRAJ4;WB#9#@AIW[AXWbR3Q&f\,16AR\S0,N?.
,8KTN\LC2M,_OX17c,,@+X\=fFJ0f.F1[2W>7#XS>9S/,_A2XC2YdS7LJX#0^dBX
a5I2^c>Q]T2MX:=6fK=cTL=1,^dG_V;aT5TK&[c[+0g_#3_4E8B23a?>dCKOP;K)
Lg]gAPDCBAY2a3AY-9Q;AcU9VOHLDI>2.-B8HW;4>V<9TB6LQKI&>K9?BG,ABFEL
MB#?W:1Pb_IP+XCd8<,4^>0>DeDa,0:[M#1Bg,Y@A\4R<H&0?Lb?_P]NUPYWTA:K
JOacV@_XVaE?Ma#YG//R18,SQ_a:g)a@DUL_7-AF1AQ:Qc+XFC9B+#_H</N1bSF(
I&[>\4[JU#.>XP0b,GfE\;JV<C:;@Tg4C-N0T2SHOgXYeW4AMg-&O.0Bf8ab0,ML
GNZ?YBIKLTLD6dC0P)CGT6<QJEU&JB29T]+D\YL1F2Xd8-][9D39.YSZKVHHD<68
(T8-F,)<GVTcCF+c(NYH@PD>0PT/]F4\^:G<_\JU4CXTgQGM9./&FfE#7aK6)N+b
0TNR-2-;=MYaE71^&0;fJ[Ac)KM.B-AO8Ae<D>#1c7:,SdgZ0/#V54OY52,;-.0b
U<:EK\FL:51B8N#?dO&G_;([=.PH=8R1],Nd&S52=25fC\&5<I1KF\0].g-6H(87
?KQ&,+]f9W_&>>6O,K+NdVDaZ6fA5SYbYbXT=@G1WZRQGbBO?VR=0S_D)9LY4BPU
HBed-3<Y5VTb7Y,2CYT]E]-eQUP04H_HCeEL(3&=BOX-PGGdcX+X2Z]KL8&LEMM_
9Ba.4e^20fB5?<GIa<V#1Id2eUN=NObAQ=Z1d+TJW8M[00N5RA=?BUTW&#;GVf1?
<-eR_7&^0^A<OGLY\D^7[FB,:3G5OJ#9=ge_4<8Z[gdeG82;ccfO1+EHTY10WHVE
5L10\[-:3fU_bKG2BSSb[dL\(ENRQ5U.=.X[Y_XUQ>S.e[0/\L8VS?&:c8L[UcUN
<(4NX22,-)WEYY^^B/YORTBdg)P\aW1Lc-P.9+F_-Fc/3;G@bfQdHGQQKOMM7;74
b]&SY6M:&AQQ(gJ:+XP?gU63ZZ(,YZ0&A2Kg6Re18?aET0SO8fcXe,Q0X<49=C^E
2Kg:eae-MXYM,d@-0+GV=&e)6]LE=V;JYETCA0RXAMd&WLOC/N(-HVL.AA;L((9M
MgX/XN7c.,+H57SQF@_PR(I-5+(R:,CM,SI4,B?R=>_TD#XPY_0b0be/cgdFZ2a0
_#bSDFLIW>2QP-eaJ(]36dg#SJQ9G#a@XV;Z(IU\>DQE+D7dV>;\^H7PD;LHSe+5
7V<R[eAB>:)MG<JIR\_3:+S4Wb02SSHGIZ=EY?\MQgHW1CMD0cgISTW>Id2R&bX:
L#=QMU)NR0cVWPVGfa8C[E;FR7b#8d)F^aObaOZEB,S4:6Mf@SN<9;P3Lg&XKZQG
5D]Nab([&L5?]=gXOcP/cJMUWf.1KFMSZY]e_/bcg6QD@HS]7T<T><2f_d#0AeV0
g.W.;ARP-ESV1QHc7E=a@5M(4#F4\0(&[)+eUO_]J1(\e#N2&cAGKc;@13SAae3,
?99dI-6\^R+LbAAdIO9N2.YQ88OLR>:WUCBLO,gc@T2<HdDZ+0]OMWT\XR?A?,4L
CFPDd@>[HF&\dgGLE^BPa4[S8IPUEI-(D?Cfa\+J=O2KFN)D8)UZB0GX55+1?8T(
1&?AA(M-UCO+7gT79\_J2Le.IIc4GB+/0AGG05.aE+P(<aC&_^7eXRC>Z+_474aW
OZV@c@B>bUVc.?@=edES+:D-AE/;JO(+#b^55AMPf4X_e)H]EPUM9E,?=3FP2A<X
B:7_QTR6#PDP#00ec?b@CN;<NfO/EZ^dUdOE?;3/,#dK6aX4G:A:+FYacXX5NZ:Q
[I.25V>LW3.I0&RXWC,3Wc6:+M=ebNEA^g/RX\LU/:6+MPQCAJ2B-6fDIG2&_N9[
7#@J)2P[E/OSd@]Sg]_G(4>D?ZY1[B@#dLG+QFSIc:QXOad?F0H=7+f-+dd3B@bQ
MN^X?89f_QV6/\0>N]+1ZH3DIf?cN@L98U0,KMacHPa)g07ed@,=5d-10EcG_/>2
OCJKAXcNGS&1<O&9aG[02PQ9>6;GE^RFD66g+?)OQ)Eb))dHa,f_,56(JO1EUO2S
CUH\K)_,PL0g(=I?+abP\b:0>5<CXJbI)/,G:VJ,e1cKd=/#Jf4B.bK]K6U#/HEJ
\_Y==ECV^De#>cF:9WT9@.8;=c>2W5NS6;FU-9JZ>PB04G5[/&(P&&1-TTQ)H>#/
,8/g&7:8JUc(J2:]+Ic&/d\)f0RZF&=E7gcFYVKa#::SP<O;eN16:NO^F-\9J/0:
AY_1@O;PZeYd\&g?X.NBPcZ?DAS#.1)U@ZeW<UJNFXNIegTZHcVc@K^1J\a.ROB?
.7LLN9VLW@J_[O<RW[B8ZV8M\-ed&&\/)@]#/5>-)@1#48>V&S8DdVF):TUb[&\.
1?1+:N&JR6-/=:08(,8SG]A\DN657S?-facfP^D8,QfeO;[\gSbfMK.ARgDf-JJ=
SaW,W3D5QRB=?]?YSUW+3#?YMbQ1U.-ac7@^2JDR?[&+J>OQbF4^=E4[9HY\^J_;
DQMdUBE[G?/OGFU9JPJ8A1;:ae1?>MS26[-LRJf5LeMd8(CfdG<bQCbf<Qf4Wg?U
A1G2g/B;=41_/DVO)YP5OX1[E-b?U6PI\<T)?C6WC<CCH3H<^2R6#XER9&_B?fK^
S,M?@Y_L@FSV_dD,:1AD&&9:_>L1<a,1aZ/33YUVE8(BJVUHM?P6Y\XW?DO2(HB(
[=@.2N[BA[B?c/MF^=I5(S8[SO:<gR^U=OI:^+?BD36)2-M.KUYE8K>@.34BX7VT
3-&gHdSG<ZE]HfH,BW<5],UF0K/50bQT8OAG]^X(Rc;[f7bYbQ-GgG/BU6=PgS[g
<SCT:EQ?BEc8B+5AED1G+@7f7.eg-:g5\JYC0]R(KS,F2G^@X(S?dBAJD]W=W7[@
V)W6A]Da-^d-4OH_901M=<EW#EcWQ6?FBZ7=:P<OceUG85(&8IB2/gX,c/e)d\<^
Z5&E1NIJPDNQVYa6Df-&=@9JU+RO1@>(<aP]2AU=UVK8J.U6;H=bF-&HF0#Z<H(/
;>/)X/-J0V?OMXBG;C^0TCeVb\9V@Z=-.dWX;O)K=+?&FS.?6VY8/.I-;HY\62ST
aT=<F;BIRKK8b7(86gARVMO/b]1T85HRa>O<,Qf2F=a8?_(dI(J5V;.TI[D(ROf@
6T-0c.T6a#0#IU7EH22N>7)-Sg?UY?_5;Qd)7Q)@eZI,#UdA1gaJWV;#N/R\@6g6
SET,YE8GOOM)10B@OX.]f6O8\,U.6;[ZgHS=>.H=(P3VX)NL5dW20KeS2b+D_Gbe
^PAI<_(b@P_VaC.IXZ>SE33:#H&3#ae)UC-.TgI63bLVKAG4Gba?1)EcNN+UJRJ:
[M(P5[8)g6;;Jg.4Q;4,9J&7MO1>ZeWEF5g0OcL@3+9XJ1XWNT<^L>TA\SQ]QN3J
PV\[J@ML->BOHO:?I1?O>E658@YPeeZ+/Fc>g)Q&N9A=+N.=cgJ6QHPMIgD(e)U,
bd=NK,0U/5AO10P4NP]2U>LdBTSFJ+eK@6^3WQH0I#eT<Cc-;XJ.07@^6bM<F&8b
0EIc3F.]9L#CTU3;-6;3f1@E3/ME@(Nb<;F51WN&4B6+)YAQ3&ZR(0&&^+^TR&F@
F)83WLQ-(b]S=G=<R3=.8MS.ec^,O;He3bPW#ALFC0e-Dg4Q>Z?1)=+bD\VJbUA^
&/Pg;4HaB7MC7-=DKE6f^35g.4XI__#SSIBVd,[S>LNb\P9G^G\NK4&GV4;MbT[E
[W_IK(C7\Id];<a.E0YI1;7GXCI8P[<V-e^c2EM7;B[)W4B=&PfS:,RD,;RM-d+G
N@/-VIK7_7L:]^^_g<X1DH2_\+P<@HFd00BKO^_HQF)X:c7gHF+Q7XX)\)ZSdc<c
(&=:^3LBUY,.Xd1C(K&F)K1-))\LJW)N;,75YX?Y7BEM?MBM>0C4QZ2[J67XE2V0
GQM;#G\.-:VPD?W_JQT6d[aXSdTd^/GMVf0LR.&2)Z5U)<]D3c75d]_RAS@BLG)L
,[g,R2AIYGK=R[C#DUT1<]-?M-E)H\Z:Z=Gd4;;H.GYfG#8^,=9;_P?d5c2<;\>D
U_eYBeQ;,J\E^_EdW0PY?XMaG[T>T6IX?K#Q/QJVNFR1VC(ZbT(2TR)/K^:6d/@>
CPg(9R3I7Gd2GLU/,ERYKP\&ffd/g.F6acE5#bPJOZ0P(-EDdA,f;T4P::^FIbYH
Sd3UFde6^3@R2QD^aIT,e]Df4#\03O01E=C2NYa&5O.2bf:bUc/b03Ea4.:._5O@
RFA+Raa>(QCDEI/,2^?9HL-5^fG5d4gaDCZ#2?.:F^SecT]JXWId:M/P^Q4UG6.(
(AQ+M\Hb+?RWgT5<A,/=:L:UBdec?-Fdf3-I.]R8Fc<b3<W.C:D@#A/EPf(Ebb.&
)7AIL[/W<fJb/(4XP[B3ga?-\c0KJ(SJY-/FR36+J3#)7W26SRc[;-TD6U=EH+Mg
g/d7?FDM,N+O>RSL;DJMWVO?^c]PNI-Pe61A+UQf8>P[\FH4:Hc_9M?>BdRF-:_O
TP[7-V7F?>J>\J4d7.=LNNK5:#;8LRGNN>2(2+C5H&.aD84=.E+>8HYWM6DB&J@)
V(NRQJJC7.B..2>#gVCfVT\F6LG^7JT9:XM])A?NdGB[WeVZR9BXG2PgIa\BV#WI
VS>d9PdA5:-#d@F(YHU&EG3LYWEN/5J?->H-(H^V.T@H\2;07+ALWdbT;3eP(Bf@
JH0ZbG/g3/KEY_\/R:bGeF8_U71Z.84aVYZU57>2NcWJARZ#),>UdM7UEAebX/Ug
5UY<ZWDfN\\#Zg[9D5b_2;.Q:C9TM.8@,?UEFXbORDcQI)c(2DJ.b0]MLCX:2f--
>2;K\,JcZ(GJM_fRZL386@71]3cH3/^YF1/ac(H.S]XXJJ-9fYS+,C+gUO+HJKM=
(DH8NM<K;036AD?4TTJ_W\-b]++Sc(0<H?^F0eOB/gX^,8_C/T683\Y?)?4PR&AY
9P_W?7L-RVBG;<0;W:)?J[fE0f&L-OLdGLOC92LVR,BP^49[38IOE<W-Q6:YYBe+
K3gIc0?Y#65_XFFCNRZX:6M8?W;b57[7.f\#&gH/FdEEZYMcLIF&[SXGNS)[05-+
2eOCYRF2FZJUJMg3:a4>S87Y]UX-_I(G2IcX?MBZVC<7_>;UeU83(2OgHYWe?WO&
;^O8:H+G1FFBKgL?Sd_FK\\d,NU+VBdN+fBXQ6W-O_Z,JagXCSAB7@3?c0,]\>C4
-(VbKIF6YS[5-d:-6,.&6_&_ZW@1_;HH6c]F3USEZ;EDA\Lb>ZIJ^7.ae71T>90J
a9,7;5G1()GC.aF/c(4[OeL5P#Z:a99I9gN6ZQLeDI/F?;g+,.O9GK+;V;g5>.K^
@?^^3_&>eD8ANc]V9cF.eZfM(LeEKU7cUHDP(9W,Y.R1L5d5L\_Z/T3KT<?JK9KK
R7_E\L9_>5)MX2+,,.ZHa(:FA:M=)QU-LB<-Q2_T/-7;5eD=_bEGMFK.U\[JJ/_H
8A@JL05UJ[?K^:QcF6JC]8AWTECC#=23;MgA#Q72^CZ^>Be8(BA5[f+/0_TWL5,B
^\dFQBegd0L,KO5&QP[HQPS.XZP<Q6@XcQH[Q6C1VK[(gEHeOBQ64dH=9VS?-g7a
H6TB0/:;O6^LD4OOZ;&](CGMDbOf19.;LDf2>0].\J7I7D?W39b[D@BW.;NGLD1E
3<+G@WFCVTJWZB#DX1H&4,D65ALA@(=B)8>NgQ88OA[f?+?.)W>8S.7\[fe;>K-;
G8MX\,4_#<JR&UMfcJ).^B.]?/)\Ofd1;a8:HBO[&/RU2)^B4UC?;_\NY>BLQL,T
_f0(-c=aRCD#Y2XDcS5LX.=F[?2XeIB9TWZ[gVKZfd_Oe/KR(:IOWCV])=b-Z2?P
X3a<DB:.Zb6I66.[eD^ONOU,PCf#QS?<4NRCOL\A^)B(ND\<SH&:IcIQ<:X.FIS@
5#d2#F0]SMC+BaO)_F,f>ReY^PNT)T#I0gHa#&7<c1-I(bXFXK&=2<4WFGC,Q&aD
K5g#W;a9^5A4eG&.g<+c))9FNVO3cOI.fT1Z>\+A#^1A5TT5:eFKOU.?KL+^DW\<
dTV;:\@ffdc\1+C-:E(RP2#-3fFYfQ=R]GJ+SVeQ+:VJ(0RAZZC,:.XS+5e>;1T<
WNNfH24gW;CP\6<+--[3&ONBUT\H\QCE\O6f>AT3S)N&W0ZCI07N]SBMMD00FP8H
2MALH&Rc#5S<:NSG99N3O#]N+VD(36NTBK=QG&)M0BT)C9Ug;7RMCV[VgO)O^J9F
+J7cb_MO82??@c?PT?XF&(-Y(^Z\H_[;93A99(@/IC=O^X>BJXYa=4LB7D@e[\^I
E&c5[A,gT]@cEBOQB>5DdT)-7AWM1c3DVF4W+Gf>eG&ZOd)>-^f?\V1.c+0^HHVS
X^HF5+M@.SB5=85J4K@ZL<>+e?EDKAI?a?,9aA>D[;:5G\E(Pd(7-BJOW+ME-dcL
XNAFD(K(2/GYQ+e2S_(RO8U967F++A?/PET/G78H]@P@/.BBY+QH^X;dT<V;EKQ7
GQ4JWTHfO?eWfIM<1EW^#2+,LIRBP+/TFY8K@92P7T=81BE&a3Dg?HF+IcB27J@8
F+f<I^-&AW.U@4U^gAJV301C86T2P#)6d:WQR5bO423.bK7:UOG<\MP.W7,B53bY
ZSGM36><<VEVE;^c,S/g;MKc,#1\E9)IN&4fQ@4#LW=a\PA4)V1^W#Y589>#V>3=
@&#XEeW?+JA@_BDW0KEHC2MO?XSSV;=:PN^2,U0?U7JCU()?9(^e^ZG+c/K+\B5Y
UW<Y4JVDBN&?8>42WN<S.V<7g8C&fcZJQ=RY;^(QSQXP+[B-L1QaVU?SIbB-3aHJ
BQD:1SS#a>7H.\MBAF>3f=;fWI-d#LL-LU[>O73@UddQJ4e18=.=LC1]9]/LG=FS
#TYH[gc@#E_&3ZSWe<0DG5[MA(90I,6JF[E;KK^]KZB&aR:dW-VTFe8RaA_[<IPQ
8[<E1K@^P7)8ACG0FUL;>?/&f^\/.S9J3=601&7#;3BYA:O;e8COZa7SS/YK/^L@
:8;D=C;/]F:&4Q5PG7695K2Lc03@=@-I;#<,N-0@bU3DWA_^W\/b]7LLMBG]e96)
M_I=&B1HEgH:Xc\:8?.JYPbLEbTOI<\2f4J4D^e-0<+,OA]L-)MIZMA^\L5:5AS@
TY2<H/GCO(C5\c=&>4)1:[KI[2<-#Rd2/7.0c89aZaA]CZPGG/UJdc,eG#(KJf16
GV06)JDg:@TP:cRCNBHa9gUNE7+)SW2A>VH>11;<_U39Q.-cYY1<>RDJ53H5RZXE
6V6;f3-ERP45=PJS)#Q\\6\IUN;([2NR6F6[LYHEg0ZdOX\E^@?I[YV-<2UDU;X=
P(ZQeS76C9/e9=C]FAYK(2:[IKHHb>e)Z.&DO_F7FA8/-9cAP9b0#@X)P3=eD]bW
G56RN<1Z?,Ke:=Wda[bH.4#O7++(GT\&N7FM?SUNLbE.-+,6g4;d,-3585H&T;Z\
92W1^dDCONUK7UE762ab.F-EfMBfSX8>#(A9#,Q75>X/Ja<UYVK.ZdU9g50fPfU2
D8(7=2KH<?[;WUJK5&a?0Rd8)&WO]a-2#LI9__&?L?@I^6MQ),HDP[)=C7ZHbM-I
N4D@Wb8BZ-(f#E_00)6\dP_2APJ_N_&RG(+OECYLfA]3)c.JED/FB^5EZR/(I6?9
_4>F:2K\=2VcS8NT.BbE9fTd.OJ][NFOSW-13d:RC=S_JeJU:PV),(e8[34&7:(4
@g6gIIFLG_BWO@+.@F:?c9O.D3e&DW/00H_QNT_B#Q.K-Y/ZMPDXEES/)b,?9F(3
RD\<QgS9NYDLZ<C8@?M?CTP6//1K9(^/-=AZBX;V,^(=76W9;BaP+gM(c_e4aR;-
W@?1[]3_a-_4dA@;-?9d7I.e9ae?/d:)9X5gB4PB<bXKPd<69C.f#\)Z5AVG6Z:O
TB^0B10W^;7X4P8>TDG=;M+UR9F\Q3MLeQN,W^93/P1]VdBYWd2)IFeGX@:RQUc,
MHV[/3A?a>V<PX8UB&-fg=T+V3A#8P55J5a(9cGV^R+H<SA4YAKT(8aXHILW7AOW
P/DZ,:C+9(?.=gIRUPfb6G;PK-S/2FO-M4J/5fBHV[BHa-_DACbJg-&G<:CbNW3[
45AeG>f[H@2^9&P,JC\T2Q@)G-^.b69UZR:H6TQ\YIJ52EUH&D^Y[]\_O:)PJgP4
Z&_,@KY7N=bTV:)E^X\FX8GaA_L.DM\M\]2aJ>E#F8X=.2?QJ0[Ng[Q=IZHI(8XX
TGe24W+M-I?(TIg+#/K.F6S^5UBBZ,(CV>9&SPPY+ZVAQK]:8F:U2_K8KMEDV5>5
KgBI4Y1(<XdPT/c-U4CcP1FJ8?7Z_A.5S]:.C;gDD;eO>09dg#+_QHEK[PK@VC[0
SD@\>QG[2RH7f_)6UQ6Pc4FW&T:S8L>Gg1XI[_aY.Nc4)HZIMYX)&W0ePRLOc;V3
UH7[fG/c1M<+5#D+X<#WX\?B@N7QL_:^VCe)+Y?T+D.NDZR/9;_^J_0e@#K0GNR/
UT0O4)IFQ40PP;B3;;EA)TZ/A1F+.H0WTY<:G,d=KTP(@b/f1@:f9+]<M:2[Sg&2
9>-E^J?b:MA-dJ[3E](PE6(fEb0<UXW]a/0AAB6L2ca0g0/2=Ha\-P(_c)#^Q+_1
;C3VU[52]]20fYG.ZJ;5HcKWfEb.g2&5eW2?PSF3LS1ZcP##(BO:>@B.(:E.R7<O
W1XFb&\T#YHJ[)cT1TJX?7F9cF6-?5JF-^QXAHWe#&D(Z_?S]]O3]a?7FQFFD##Y
KR\?b+1+BFRSf:C]8O..CR+.HXY8T\\g6M<E+50d,g(C3?B[=W<A.>)QZT0CT^PV
S0@ED#N^B2L(=M>4LdG7&+6/Z0O1>U9Y=>CM[8O9Z,RM5R=<aIe0OQ?]He+c>c@F
R1@4M=/_YJg0_=[b+K3&[[\5cEH_fX\VLEVD7FSVf27b;QH]9A[9.PSEc?Gc(OdM
O[<aNDDc?3XgIIBNY1;IEN/H?6FBa@X=LAFL?-?N?A#(&eGeL-WB.-18fKbWR1;\
]]:>>1g)PXeg[KCD[ID#([I>V1U#_bV3aN-3UZ=[T&VZbeM/^TXEO4).?Q[?,SMg
/0.B-[TKd=YKMS7ZcM,3A2b0[Dg5_0Z7Y,7&.=UY94S.Ja6&Z3<OS(d3RV&#I4OL
4<(4K1ZEdU=5^WT^3(L(7aeON)Q(G\P\&FCU@O,?M\0YH:T2Z)#b1PP1IcB7X_KO
,[@C#>O+9O5(:W,?\TNQB6C#E&,4WQQ?/7]dXDB30Q;eZ8=W#[8=C)PP(TP1cdUV
1N0a3M:/V.R][OA[881>;\4_W4TA8.bF/IcC@;4:.FB8W.3(MXEF=B.;<S4CY@D.
I+UM@S2\aD0=(:J#=D@[]gTg[#_eVPgC_>+(3[D]<><Z>37\;[8QAQWdKAQOSd^>
c#>O,Cg]AR8.9a;gI@aKX2<12-G)V<aEU3PU07&gLL1JP^#4]80F@M\8=OL62fQZ
+BXeK376JNPNJJ7#E?T\K44/Ra4C6c]SN[R0g0PK4\Y\7+9Bb26X;L2L7471@,\P
[2:FKAZAA3bg#0gRC=I11HM,615Qe&S43@[R[_V;aUFEaYgReWFE1d8WQKPU=YZ#
(;C79\KaV9;O[]4&9IR3HZ07X57>f__EMX)/VD#2gC8<R3KR/Z++NUN_cOgL_417
9/>@PcQ&.0G_1GP^b)R)[=>BF:L>:=CGc[QRSMN^dg;\ae96Jb,4:]La58F.:7V1
7+Z6D3:QOHIK?fL([\#cD-?RRQYG3g.+TH0I?a?X6^;^d(,8L^B=eS4+UXF7A2#6
7B9EA5V0E;\>M,ITXO(b)MKb:X]5-<HI\[<eX1gOO(LdT2_.OZHKO)WRgW(eU_2c
afD&XFbEAZ74NPD+^)YgO4M,bKK^A^68[,]:K/_@>a<BN^)4IUKc4Q.G2S5^#M+)
eDUHLFX&@6437M@[8>S\L^::PbZ.]SB#./gc;,E@_EY];&;6&XdDE_DH2gdbN+@U
:3P#3?[@NV[D66/WO]_5T)B.55&MUG(^e74L#JC?LWR<IW=Sc2]ZO&U,g&9c-(9)
-3IGCP<@95OSJ0D@(METI/(gM41PW8EFcY1bE3LfF61VM3M>=bS_Dc#-EPWEAN]V
DL/[I=2V1_EC5Z-+S5>XfPbD3Z1R,JW+OWARO(VV?P2K1MPe;HZR<H3Z)=CDOZT6
@)4HQDHB5]>H0YZL3VX9_5S;#[5FISXZ5f2@\CSO6E/W@N;O3I@R<O:C9([LWYUe
H8ANODRXF<(=NH(<<GX89?=^dg-Qc[:5U-e149_(,Q[6Z]9>1e.5gOf0Y?G&^T[K
GcE=.A&4RL#UDcA8Q&[N9_Jb95O1gB9gS]/P2YZZWJ34K<IQf[/-E.4,Z/CG3R,&
+0e4]GL<7,X]09c[RJ-2TWN:c=[P8RBBdLcD:DM1YSIf=C.RRN@R_gHK4BZAZ&V4
YR<#0R(6JAFX+TNJ6#BDB>,D^;eHXC1(D8-KR\HS3;5Y0\51O@4&N;^HUBD6Q6Q+
3c)4fU4H+MPD4[#]e24daU;ZG1&Bf9UPS@O&K:T7E\&/20g^G#0Nd9?ALU^#+6bD
SFA6H]WVL@PbUER0cfJd>EJJ@U9M&@.8FKZ?MW/08=5/RBGK.#VP3P/GC#Z45YA\
&SP&/^cENK/H\IV<117?9UK_)8e(C:=4ODQ.>N2;dBdUE,aYLZ&Q&.7W:?gI-,<F
^)I0L,./]ZH<^RZU;S#UMFOXYSZNe.8+;[R[Tbb\/fVYCL7=#dS1QK^VI\,A^3Q\
AMWOa4L_-8W<gN3\AIM6@FQA6<d[IcJ##^D<XbD5Vf/E6e_]gC&e@,U&UVS)S;JK
E8#BAVNa]&/)8JY.+9R\&G(W3.>d7;7PC4.F,5IgE;e_ffART_?F<H=?)S4dR;VS
=c>.M2>;MU\EKGd\g4Q8MS7C((=\Y+J?X056Y=EJF]3JVYE#(=]U#S6K7+<+&FVY
2Y33/7O40OSO2G@?8U#=-f5X?((77bPU93</Y,HKYS9b>a]R72WR@cN2@fF_7FB\
SUR_[ZS;<8?eC0Sa=5M^dPAJ#KHMY;.O9f0gW#b]N+\5@fBaVI6>P[L6@dG:?K)B
^LaM<78GgC&>fV8D/F15H-J+HeI2YO:]W\S8NPVGOATQYNI?,X6>^^;.GZPE/@(\
]Z;FdK<>/LI7Q(9<VAMN5FgfV253-Dc0Y123H31B_0VFPW[&eO&8+_OSCCMLEYI4
eH]TQHP+7//(+/[92bC[0K>WI1R,E,\).SZgX=@,#,J\+4&eLYc1+G[B9KLVeX;N
<IF83T5+35[HS-4^B[dPeKC4E<I<KCOIE@P@AgOe9-7<_&3C7FNJ-V4bJD^/Tg;G
G\Wd99_B?fNNg1RLS\eQCBI4-^UQ(J/L>Lc0d9CBA],B^)4ORKaX4DM)[GF;3U\\
@36B0?;,@3S8>1029e0,ATYc\@N_g\(HFXb<Tb8=J8D&7^U2g5UAMM>gO+:CK_bC
^fWG@F5<XYR4I1?AM<SOMP[7N69f_]9-U6JG\V,67>T<==)=M@//\H14d_/+X?K1
8YOA3SF7AMQ-U8H8g5Y5CI0<I1_RVf8RIG5CPLc39DHGFUD6Cg,&7]C[d28,P=C,
+-O@W7/F4TJ=W&9-L2(?g4Z&PeTQ)55>2#H74J\=8>f0RA9/J8B7CY>SWaF;YKGg
_S5b49X8M)dAHffZ<a/I+/82a@B934UZ;6Z@Vc^J/G7I<2M>]f1SD>3H=R6M@Vd=
<(70e6+,ZgSFMQS\09G;GW9&aG0f?B;\F4/[(]Q#;P2Bd;4)7@aHFD.P7=VbS3&0
A9_^2(4&0,(g8OO^bFH#Ab)K/VCe,ZKMXY(05^6BMVY5F8]0(4abA25BSBT(GV&g
edU<Adg>cNH[TKV7f]cAE1,J<G\TL<><)P42A0GXb6>++3),2D+TO9J.=b9,Z;T9
d6W:&ELCaa&]>CXg-/U1]c,N].bfe:f]BC.@._7;Hfe12bY;JaW_A:[H\ZF4ODJ=
-@@e3,46.\5c39ICa-SXS(7LUL\K3N_4[2HAUD2RU>8;VeFGb>Y9bD.TGW-[&/Ee
OOaP[Z9N#@OWcff/De;K8C<HA@X8[US9@WX:aL7a7a44MOO3#2L\:3\(eY.8M3D4
,[35\ZLBO],87(U-:]b\.R?.HSCT<4/bF(;EU+R>b[[5(8EE:N6[A&DL0GX\<1TZ
J3AWH@K_Qf/(e2I>^a28M;UZSJ](e;5=cD(NT1BR?)2DUR9NG(I\-@#/-:PV-0B5
J0<A[EQ.9T9A7J:HaG;,CY,=B#2E4f,-A_[F&L)-VM/>3e5R-1+cC&Db9RT5PQQ;
(S[Q,ERA5ZYg_M]H,+4[)-/,/E7@?T.E,MOG92af6+-&F4M]OUU?Q][IW=.V@ZYT
)K8&/77C)0\31S,8c:GYE_YPJ4KEC1XY.]>1-#f9?J39?cRgY]?+EWB73d\Y?=&;
8JA0GCZ7Qb#[\J@_/[3C5.DTY^\bZINcYcT).UQP08f=9e@Gef<e?0?:ff9dR#f5
N8ZO6NbR8fB49VXJ;/-X=[=K8FH0(#IBVfD.?Pf:@</:/K\T[1d?]^Y:1/7\b&QQ
3Z_K@<\]1A]&Zb(IU:g6?OJ/37g/)Bf,NdR+/g)bZ7b@Nc1^NI2P0TY(cPb,-AZ^
6-f,?3.PL<Ig/U?5gASBW&b,[#cTS3CI:X.?A8:(9fgTZ6:<(eW:^1HJJ<cAdGHC
(c?]GB9=?H-&[P^/15[gEM>Q@Y=VdUId]HOYA&8>^1,GX5T&C3Jf)KCHc0=1<:[b
cS[^a7YUVGGXKRTN9@3_?bBa)B+\dP9;N8_5<XL&GN&1H;E2TDUe3O^]6a>Q-:A:
fRVc,b;Z([HK1UQ^cWRY42ERS>^C[)K+ReOET_c_K1W>Vd#0f#N^(L.CRR&\;&>B
VbP=3RJYN3KT+KEgMW]D&YWLe29d_<IU5>CBCKSS44^_=UN::eQH=Q5a[,V2X:Ib
U,g_WG3eG(3Ob0]6?dYX4,>0,5fWP1_c_(+WU+aI<f-1gQ6LY#2:WOIdFg?_(M74
TgJaf^4O9MTTB;0R0fKI)3MebVT>>Jf4Bg:9X5Zc.K)1Q3T[?9Z1_\MV1E->aWAH
I;f4G-J\f/0,M#ZLQZK_5C9?;bbaJX_5_G)JR1@<CdU2KKMIAU<8+d5Z+NaQ<Ad6
Q81KWE[#/E.Z]),b6U5[eR\(HO,:A1<>c]KO+FV#gd:&OY1:D8AK3\NOb;3.dUD2
/O6DPIYM2Uf5]<P-D/G@(Y]b1P?VG=c/g(3XEJeg37OXE>H;-VOQ6YNAf5=+.f<B
<4D3Zf)1f]df66O?F],F&@DUI7bL9YS^BV?39(^4+DE7b[5YfQ\f4e7e7H^>Z+YW
XIfI??Z[@bGGCQZ@,SeUII&)1,Q^]/+0e49J]-C1@CHLfN)4QB1fOH:e-LAQgO:,
>TZbPQ^d.B@cS=cR.L;U@4[(d>/[5B[HQ..O2]7-4:=\<N_I1J,Jg/BFgHX@eBB0
aUE^4(=_7-7OB,Z/<.F+3Na]>>QN+AM>d;(ZH=/G(aO3#.g&bXe<&b.3Qe-\+]PE
Y+)Q>2]8=e-=KP-,fe?M9agFg]d,/G=4/2LF3&\<NYfX]AP(LOXB[WUHG&Z^HL&+
a\0#S3@NF3CXK.0gY4X):Y:CD=\EMS<T;/SfIMEd\-,e.f\@CE\5/+T2GJ;RfS^7
HLEXZ1/?_a8S6ODcGHf(43^\YcYGg;IZQ[-6,WBd@.P_VWK.V.;?ZS5I)b.21:&R
9U;Acg1d#YgDP/P,3[P[FGPEP8JURN>^)))VcG\Xga\\8@VKeFW[,O)7D72M_+JP
]<e=e(PL5IDNR8R1_YJ?K68D-/@FOD&Q?@15]a5^SS7GCN1NQ:G6aI5Qcb-B)eU?
CKT..M4C/72gK?aF<b4WFH8ES90b&8c4f[&W7<ZK)<IH(Ag(#G.0&5f)TRF53Seg
\_R]FT:#VO=)@g>;&?)7;Af2OYV6M.Zc3V4&.I<^X1\4.3Y]XGdZD(6JZ_[IA;Af
H\O,HYL75R\:TH3f&;I3P3PgEW2c;\(LAIa;G4I847>_KCf@#(P#YXC9K[V4O@:c
ga^UMQF9+^\63f.a=Se5BM<HU-Sc^OBdMZ)JF:KNdKKZe1&aWQ=HaLB;-=]Rg\X9
#;PG&TeP<=7NK@-BUbX@A;S]202aD5=f(FB1gZIT7]F6VW6F=Q^B+U2<c.8R_HAg
<bA)N.W^4HHML-\R?<aDbb,bK?JM@)<>QcP.:BD#PUV<:,^-:_>=][&g,<gIfE:H
Z(:B,-@++];f386HcbJ,J^9<H:;f<[PdVgPKCQ3bA&^)M@:g:RN_a#&G#a2PaZ<.
^8XT-)f>O8O[A9#W]<UT1;?#KL1AYIQg@JVP,KU2TB)QAO[E#]GgcJ?>7/M-:O]H
a+2=>)&2\.UY],@;U;a9008[ZeW5L&1DE(cf-V,BDY+G3/K\UZ/N)76A45.(P\#+
#L70+:OReACU1OA?cXf<Tg5eR;;^[L(4+f4]N-DD=NDKf<[=6QL_<5eU6gfSf6EG
W>E?J;Q=EaWTPE1>).2?.6_;6\cR6fJ0W&5I1>+_U@X?I;<U@.X.-4cDg=9SGS4W
bT.a3AgY]YD(2+3FHKg2J.D,SN-e9fF<<b;;c?HFaDBS&eQgIf?8Ec+F\fD232aK
SdJ&gI)B726@=2/Ha24:H8-P7fU@-#_Df).@16<9gdF,QAG^3&<c.V7)gA#ZG>+U
[^@[B4@e_8gbB7dAZg5R\KOQ339+-XJM?78[GZ#-J3_HUT-DFSZUM<>^#GO^W@4,
9,;^BQ0->^dFG)?G:-VD1\C8>@MD/#bVKb2QWgg0BO#WEg89]3@8bJ5>_aKeN-4X
c>-EbeNfV0gW)DMT^b7C5Tb#.6^EEf/15J<?b,T>J)cfUAPUQNO+1D?MRF/ERULc
+YF0RMJ#):\<:5DBCdS^H]6R8HD-FXY@(0XDMQ9723e?/PR.XU0JC2VEVB8/^0Pb
]7B,&Q)fc7NLT8T)>bf;D8R->HU\Mg=ITE_>_2dO.(5&5=W3C]#gVZG@CH;I8WJ=
N0F),/Z]cL[\6BJJBUA_Y[9;edQg;<-29V-+\EJ9UYFXW9P0H^.)B0;QY]@M,^d[
3.2XO-\<TbcA]W;NR3HLG-QF;C#fXe@CI87@b;Q2?W7T)FV[f7UfHd7:.#FZ(BA>
[5CG9aDMZ^HDCeG^#0V_K:V\eRBO?(@G9QQHN=;,?3L.2LBLQcf3/EX58+RM7@V>
GUJ]\A)REKcC-d9Y2JAKCYT9)]8EQ]I[4a/>O^KEg8K1B814TFFUNWTHJ[:?FGP3
:D2&Ya,=#C(@<Ua]6GZSX==.GY<0^,Z7@-L+:M=BK)T?\+K,]S??=_R\YWI/D&(d
)^SW-1SKUZ_Wb2_39>FSg;N?f:+60@9ZG\R1#GX-IH4\51H>a^Y@(e:FR;Q:[RD[
;NPV<bc(:Y3;]:VS2D<CN6Q#&(;<\UA9QA;W_4gZV[<U+AYQ)B;_IO3@_-R0I6R(
ZI8ES@WF/=NM9Y;RfUf.aJQ\[@DRVA2(Dce12[=-L;QPae0EF/8S>^&2;-FEIM/?
6cVMK3M0]CTIcXHI,0W@>Jag2gNZ&=eUI[;KL9/;UH5\YFfM66WANN>HQeY1-(ML
R&,&_K6)KUfg;3Lg=]dfL)864d@S(de11]]P3;aIX5^a-MGIgY:\#O&3AJ@ACdDJ
ZdAfe0KI;01JX_e[I7Y@A<.W@IO]&7((fO:148PTZK6S:gKP)OaVHGWR@f-L9I4G
HZ9NA8a@fGACTHD2EUL;SP5-SO.CUJ5,].Gc?XZRab:[7DM9&2_QG,+?;2@a#L&G
M)AU</O#6b(Z-F@G+Cb/]e[g&)3Z-1YN)AdHZdQ5MJ-)UQ)<<A140.,T.BBW?)d/
:aY;>AT&ACJ#?G9],OSGXFb;Zg/C;VdBVRBC@^#d301>#(\:c?K#3G+2ECCKK.PU
#?dD.U&RF2MWWbFbK(8,\3:.?6Y:Oa8_f2T?SBEe024))L^[c;LR1/:8:<G]QeRX
a+6J?@9Y__F5@DLFLc:g2Cff=cEA75fe--0&YM^8@8ba;,4Bd8^1ebD)+XDDSDg;
C@4N-,WT\J0@7;VT.B.0-ONUb[UHV37^QX#GK6fg?RPOT-\M+J^=dJf_&45M/(R6
8>8<MQV[N=7VI[ZZ6b5OY6X)40#NLQM0+IYS4^HBH7Ed=9W6FfFQTe)b3=/(EU<[
Yb.&NNcc@R7/gL0bV?+H#+aE?>O4TO;>^07-/ecOD[d\[CE[OK#?<ENE0[^Yd>CP
dM:&0TIH-,D5=ENWJT]D4O=Xe.\1GbIOJT](6TP:))M6OL+C6bM?U&5Vb;7ggXS#
BGH:>1V=f^S+6a#[2R56ffgb/gb3L44e))RT4\G-K@Ef8HP:_\I_G:?C<(0\8Z)6
LIGC&cHN]5[[6K&_e3TLAHPQGTF348\Xe3E+PEY26\14.#Z>36f@^;1e@;]JP[&F
<Td;;N(FT+T=#1GYcC3>J[ZAYKV;4Q]L_EEENEFCU#,F#2/eQg^L/b?O^2O:gMfF
MLZ5Z7W:dP:9],XJC3:+Q3\6VD;D8eSYD)U^5)1._8Kbf-D-(>?aaMXH#g9JVL-g
:]Q@f/,QWRQd\ONV.H&,c-G<O-FZ3,D0)++Q(R69.(I7S5X>06@d6LO+;O3/5-6N
e<&57bc\9C.>(POT[P\N3E0Z9S#BYA[F^Y&(&Ja]LM=d>K3KDWc4e#f[T_U\(g=P
AH/c\T)+JeT-0b_R;7J+D^X119X?:QI_M8<AB6/,.X2(UCNfBEd12KA7;];=+]XH
3GEYffR:f[cU_/b(/Q<#:0K+(N,TU\gbM&Ud/:B(#YM?g\G=Q6LfWFO+2G?Z3\ge
CEC3X\UUQeLP@O3)A3NA^[+;9L4WS+#>5KX=0&7^-;fTM7\QC;e^;7eZKe6aL:TH
Z9;#^=NO>Y7aaQ&FW.AE>=VRQ2&L5IK3KP1a6G.D]IAEN5C7-.b&/HIJ]@]g(,Jg
M0.SULR;6;#HPIeD6==R8N?5_bS+.JM&V3#<9J&UaR0gE.3-QX9)+,F?;&_KCWL,
cSY7F6gcGVD,A;8B74dVBZ<U#B3R)>_QAWWWd>ecG=O&2=O4a6E8J>.RRSU>CL0G
_=\#Y&S::+bE8JWc#-WK:PH\8)L,P9:0T)\M2L:L6)<2M&\1#.g#ZIH=LCPVX&g7
g91,c=7P)9>5:]K-A\9L=K6^459eYFB9K0a_g/+R6):_&VbB3^>FVRW2Z?]_Bb8U
BPaJVf9)fMEH&MX:DF6R4V]Y0X<#\5JUD(&.V=e>NS_Y@M5/D<;R(?HMRYa<O9N5
/]b2C9EUZ)=R1Q7bFBKg;KUSXI@A&T0N;b);+-0a^^Fe&9#Y)V/KBO)H@N?+^ZM0
R5.(Cc]Ad7-b?25V,YU9/L?HDb68b?]=G0Q#A3(,VR+5\:Y#VeJ_\Z9M<O&08bd/
;ATeTUg;OVBYR?>X:]R9g.#JG1_eWR?#-+SK0GX6ZgRGU4UA)ZaK^E7?UB\>C(>D
P[3OD>eJBE55R#7Q(T\6)/?e8.J<+FAa3L[J_5P7UF6@?/^];R:c(R4GadegR:GT
2=7Id[<.]GdE2NgV;T=8K3<F(Pge,NQ&37<4OEaa5H<K\<:f7NaM)MZOc;7^]FTB
HgFf27@(2J/70Nf;1=DKJ.U[8@8OO]ccLS+7S_3VI_8SS5I/D@6CMKM9H0IdQg(/
42NB6?<=7>,O@G?CDG(-2;g/8]0#\/&ESU.AXEc4MMC&Y/\V.R4Z@Bb+Re<X,G5S
Q=cSK#5\^<QBdB.@+SHCLP=:4GH,MKOP@WANADGQLYW(=KFPO:2WbL@8JCRJ[,a(
ZNcTcF.B<b?\V8JB9MF:OB>:4]Ca4+He3Je7W4,0&a))A50,]=WZ7\_feZ8\V<UJ
DTMX=c^c,5QaV]<b9H61PW@DO@\2Rf4F@SF_b]I(L)PSN/^K:,ZN8XC=@+S/JO&)
9:,&)UH\Dg;.d5C<.#@1SYUBYP__[9gEPc//;QFcaKI7>XK?UF#aC_NcG89XWU_M
5JD9SY5C03R)>AUAU62C.+fO^HLa=,3JGO10e6.H\e=^Z?5AVBFPf929a#c_.Q)(
7.gQR>5WS.c^]#V0Y[IF#NI\Y^M4KfDP+-PE.[[Z_,;CgL2)1@.fB8A2?04YJ=;7
9&fU:Y/AD^G7_L^T=>:>(gCVYf).W04KfSaG_0WZIeLN1CUL4O:@7^d=7G?DYe]4
6Zg>_@-WZ_,#HD&fS?,P&eT@(U0N+PaL15?R7#V7G1D?_3J2.LM@5&=ZL3/AHAF-
?d:MZCd\d^cB5B&I6P[gVd#e#4LF@Uab,^[AW]J+e=?e9Hgd9;XR1V#DO.3(S-7U
gJ<D3;&L3#(9<EP+\QGbE0d)QWK3-SYK&Jd\Z)0EGVDfG#YQS6;&fS_R?Xb[(A[T
[_]8#M^2^#@ZAEMbH,SZWHZ&E.g<gJQWYV?\USQ37WS5G#H-R6].Q.Jb1=Z.f^]B
^M]X3g(:4.PPbB^GVFZ/I->GHNG5I=H90gbf^N_cI6aH3aQ1Kf;A9>Z&#_2\/IDe
U=F3.3A,GX7SgIG;c-]Wa^J[+A@\-bCV(S^-BIWXTMfK81ML\24aeg5g<=.W.a+C
&SYW4_-63]EUP0_gD+&cU[F<>Q,B(XIYU,ICP((C_>CcU8-H#>9ZDR/1DL.+C_0U
eZ]3M+#I9MW,_L6d:gCKX7,<<f=C&,SO9:0;QaaS)f/[<e8.,G-/+O&LLf#00K])
fEB_dWDbbeSB_S)&[9(MLeXbSF);&=:&)c>P6B3YLRBE>[S6V7g6<9#RNUQ40PBK
#M:NRg=S)DfeA.DDHa]#e[6-G#I=&IW.KKUXM++^<&.)@ReRH3(ADD5UL?3_@BOe
&@=KB8X)g@Q#]PB.&aYV#8a_13PW?D4aU7U;Y,<I^BQ7)8@M=.Vd=d@F7(6/>Sb#
a#6GeC7)@.A+)B4ZJQOc&.CQF\>TJdR-&-De+(MD@fUWD<e[[_HD<IAT(((RUX0U
MKYgVTMMF.+0ffHJG-09>FK-R@TE52223c:?16[?EaKS,V/L?:#E4;-.Gb1+D&4H
8cVA,GSTfQD;d(PBB=7=#N:-HL>cG8C\4Ac]J/Ve(KQ6Wb(b>#f;<09-ZKBKMJL.
McSBS;/=FC\5:ZaBH,+&W;J<=RgP=FcAg7YgJgg#[eVTEUDJ+3;?#:Sf</eLF83K
,B<J()6I#P1;9F1b;0#S&A#V@Xc57KC)0BNU5Fe?9GN)@FF6FH0;0)KV0DB]:)9S
P)VeN:-:N/bFU6E1Bc:H?eNe.G=(_6&5QgL7cW[\F5(b,/W[Gc[I-b&Z.DPDQ@eJ
S>9;+^0O.V4IfV<5[[I(H2IM_PB,N#HS(?:JCVcAUcJ4]+\4,Cb7fWTV@PV(.:dG
_Q@#A_g]>[0eIL6DQH#D8DfEAEU^:,&Xa45cG0egIe]_-Gb9bb&JG[EZdV8RPDE)
OWR<YHID6/DX2I.SF+KX855g248XK:c[9\/?WRZAAO9F.-;a38g\d,_;Qg@(/GfS
5SN_:7IPW+6NG<]E/-YN+EJdB?Y;LP/>4QS-<X(,9(6@HX>,CSX><(1RX0#XG1e7
cQTTdA#db0A4G5]R[P\?>E7M,F(PZ;=2.ac71VWQ)@2C?eQ[OSL#MN2ZGI#bXHQ5
ZE>UPM]>-TffQT=>-_=,fCP)bGY4dB]W^0c\@4WcAJ3a9\N./_QAW+H=,\D0W3fJ
a@U=PFCWJ+5B&VE7H,E085[R3V,HU5^Ec@L1?aPRFQHDYKKVX0;(NPJf@DIP2AaG
\9&FJY_\AIH+#KON.g43=g@XQf-(XDVafSVL_@]9X1:#KgL((TO-U.56/C):GG?K
d#>8_+,fI/F[aV[Sg9)g.5DDSU,Q0P=a@Q@.EgV5,ZAdP^Z<)\ce7BC11ZR:;Sb&
84N80&/bd1<D3654+CH:,5N)G?TMZ7,8cdHB^Jde1dV6[Xd\<EcELD(NWBTcF\PB
W2[\S[;[b?3R-U<W:(,00HF4aI:EVc6]:\3:)fA]c3:c&(6(.,POCRMJGVG,eGXa
edd()_DJ:X3CR+aM&:.C9?&-[0.a0Z@GM6:&63b\T.J8d1?=L8;Q#HE1B,OO;&JU
Ig2,cS,AC4\aPV.?g.1TMMfO6FKT>DdY>f;GcX&U10Y.#3:&D5@/I+T^_8:9V8Y?
A_SadX7/</(c>QMLOT2Pf<PXHM6,&KAWM1Q=3J89IbWgWdMC@_(4GAH\EQP)^B\>
?Y&T4PZRTJ;2b<9#SP5SPI?W[KD-aMBCQIEAe=SQ)EJaR4f6a49fS\]76QU7VW6Z
9(02X<0\.#4.M0):KMJ<(8d96YLVaJK8S3322Y#OM.7bALb6O<;G_J@OUR,&RRQ:
K4KLN(1#:)g\HXg>,gJ,7&L?f6FIS8g9DK,U+]gFOYFg--+g6>8)3O/-@WNUXTaf
b3YBJIWH,29#C:&b^83,9Vf67>:JQ?#;N8YEM/#DBaY6]Hf/M,,H4QM>I)eJ7?g\
(OG6/RK9)HDBBL>faAeD7^[eZ(O-Kf1Sb=RIa/WDBHgAM7J0G.U:8&7(12g/C:Y-
Yd#A>OCF)_IWJHG?O9bJQUT?-S<2a39;Y\d/T#W\]fKHbZ^]R2X2DD>f?MFS#g8U
V_eA\]R]@Z??,UO7#:[eg6.0g-H6(:X-W92fgZC7fG,Vc0gc66HWE84&18C6dQ:b
U0^-E-Y]5B<c<gC\;YIW/A8^P]JHEJTO3bc(.)BURM-SR^T/9A3L7O4FMMH<KQIQ
]T)@<6[5)B=FJ7[TGG^b)gRfOdE]SCX-,JTM(/bdO\M^0)F(#a#:9a[gM<H-[=D,
=M/Y/Z_K[M5R#fUWa5OQ;^2.DFNX5GHTOUg;ca_30R?0:g)MZe[gA?D4@;6d/CN&
Qf_EKIDU>;DffY_2Me@HG[]^0NP1SdQDNVbc?&OHB^Ed.7eHS;J(]TUV_eM392S2
P-ZV5(X;2V^7ZG.[ET8BeE-&:).YC7Q2Y)@/E=<.[-^/b=;,RKQ]4JG#@,UVMQIP
C(JX3aY([K@/&+d3]5@9?F8,He]EHH&W0=(WPC.8&=+M7MV>=)Z)OeCVb)57ACW,
&=c[UK89]7@M3_YSRcZR<N,4gg_N5f)aMJ>Q7M2T)4OMTM<d59^D\bSc&LaINU56
d]Ae,CCT)M3@&dS-MOXe,[gGdf+Qb1&+aCScEN7<d6/QHM&,g?8)SS5^GVP_9Lg)
=[FOJ=5fe>9dS)+[5SCDJ)F2X<\#]-gO_\QS.A/@[/ef:AgJ/]+MFXdU1B343Wa&
7SLE:,e0P@V@9B\>HNHNZ.JXVB@aUE_0KB2V,-Q(HSRIdc2LRDIN\ga5c08Te#9X
-f\Da+0-.HOJcK+JIIWO0Mb)9[;2@YCf(,C7:8GRUSI2:6gP.bb-)Ca5Hd<b_Q&N
aY^8GGL3<EI\O]@bOcKdeNZ;D\9T\&S2;?-eb5G2A9Yde7AU\3QIG=PDD.fXI6<6
R:5b551TNFF/AATZIV>\@KCIU#QBS_9CNXd:F0JH((aF3aM&VfG9d&7a/V+IDI:(
;V+F\+@-@#&1f?F&I.)UX_g5@A2MVKPb\0O8;RM+g7RL85FV]?CWd0S.b\GdI8GG
SWZbDWJEI?])T+,g&=WY/gJ5-Q:?M\dCCbaE)@1W/5_5D0&QM2MK_.e,=gDd](eb
.Ua6[V4cJ-BJ5N9639D?ZHI.f)BAEA>@>W];Z5PD>]+ONV[U^Re&Af))Xe/#&1(#
TB=G(0FM9FKD3GN+X_/2;)FWL7K;LA-dMHC_=84(PG5:45\6\.8ZVg?5(a#IM0C<
7/N7cgd#<0<I/TZ=5QNf(4):bA.Sf#)=c)A.M5g]a9)+f[?Z\0S1TN\+43(;>EFG
-f,V.0E[@:JO;&TCE16eT:)PbI3F17F<Z=IZ<T?K@Ra^E<56J)[1MB:?&0T:9DT8
18VCHd(Q,<OT&^,R9>K5[Y/c#;R7SY56_/G5=g<cRb:JYPVTd_Nc@>RK9U@O7LAX
\F[1SgH1P+GECZgaS4N]S71ESHHD^W3;F@<QDXDgH-#AG69J5P^MKUG]4Y5,2b7b
C_^)@D+P)QUB=V6H5DA0DceI:-I^Ob?70^O35:0<Y3-IB(QY-0e(G=Y=37;[[E(M
/Q]?)cF1]dT2-_4;/NJT>#(0;f#XJ+;88Sb19\QeCKEO_>5gKTfDZDKYX[KH2N4@
X&aVB(CPFU3[M9Q.0L]Wa1NPE=NT2#K5.F<+Ca?1E+3W/c:b&LF9(g1gg#aPK^TD
&&aNX&]ecRW?SS_EAbD&L#-3/F3@AF\HcXM)-@5?QK8Q-0SWMT><:eC9^->]6:,4
6<W7NHBJ9>>cA?G8C+TKF^c\)bM,OFVT7ce:d-1E3e8WY;(_J3A2U4CX9SLIC]/C
&Kd\e?d<XZMg0QbcYA(6\d)RMD)KZX&+B2Q9-JdG.SHY4];5b,\,K3/7X+gS41FQ
@[[&,6[<V;2]OH=8<8a:b0W\ZH[7P,]e./]dB=HZW/>ca7PI8IYTWUg\+4=L<Y=^
^NORcfa\:F..Lc.@B5YVc,UD2\K0eUWWRcc.RH<f<T]fHQ_)HY&E/.#EgdICD_)Y
/Vf1T_^:N(>92:<?RI]G^PMB3\X0^Q_T+9G80VYfZ:]_RE_D?HY1#G\E3bd.Z^O-
Lg([Y95AgJ-6^\CH-W3Fe)&Q9B+DdQM_?f/8H)W_54\dHI_7>1ZKDg?OPgYdBR[<
c&f>^O)QDOIe(5QFVe2()X.d#PBFa<eEB&F_)S+[:)BU)gWd+KZ:L#_Zg6c81P.&
D<d/<8&Z?(W^(f0,cKEYO]Q6S3DVLBf]D:5OKXD\2_4X0IG)c6LYO4R;XZ]HKTR?
KD.Y)E5Q(_>0)?17(DCCW#P]3L0K/-XD6]NLQM>T@1cW_57G4cT.3C:fd:9\-RD_
WL28;OdBG>5e+-c;V6<GB0:UQPOXf#7G\]=W8_RaF(,c.2dbG/KXa,=.Kc8+G?#.
E(2#XBJ9>>;Q_+BTC.>#=XS4Ga#HWBcWeT@cAAJ^&X4F7EFcU)DG9#L4JL7M4eNX
fGZg&MB[fG_15Md]K&gaDZG#I)6I@47Lf=.Dc&_2[]AU5gOUUUOB@de55WY7-^Tc
dG:_OIgA5K]6Mef-C]gCGeZ3,CIJ//FfQ>WId=Ae11<1W\SI1Sfe<W?C(DebK>]I
aK)b;XdD7_40LBNIcP3b7F]@&+8:7ALJ._BA2+)Z5:2_CNNG0bINaL;]D][T3VV=
#:5++f7Ye72;9\KVbDcV4X[W2Z)O2_bPBY.R,[,_82YP[J3IVG-F5fYb1g#A4?eG
W04M?RO80D=d1H@TQU>;QIH@EKdNFe&YAEZI6.g@(AMFX=&>^bC,K0W_P:EB>#@1
EJM+Q.-F.@6D<\<256+&T2UbST?S]ZVO^d=>9(24a5GL..fc>@J#\A/N]P,=Z7e0
LS;.Pe.4Q2^bQ0C#1@=((;K)IAeY?L1gZD48?E@4HP@NF(<MFW?EKZ+b^O-T(e6S
-gC[01/W9C(f61[Z0GT4N4.F/=1I<]UAXGO(:BC;&LVRB,NO<S><gNJ(UJRZY^,G
17):Ua2?B-@33XIEe3WOG)@M(F6MA8+TI7#,)E49G+J]+J^#UBLg=-;QAZN\2d8/
bD3N&M^fK+CZe8Ae:K>-Sdc:XG#(aScTdB8#JaF,N\ZP&H#cfXPNMA5,HE9&dbO5
-V2I+XY1MHQ4OKI&XU4<g_R[<^Ab[K9E7gO0-=Q;MWVLVRG69=NeLFe,M#IU7FAU
35\VOO_R&@,d2-^7]Y2:S)a>eC4Wd+a=#fTgf&P1U#L&.aDe6&]CSPPg4X(>W(cU
F5@#J-R;2NNAWI6(Y(8TJG_G=cdO/dSX:eL[Sa64;:[Ke^+OCI)8-JfJP)^SVCCV
<>OV80]HfZQ=-.WN]E81GE^G=5bCQL1(</#-Y;5NH9KdT=#RS]fUGCP\?dZ4)@RN
+D2b@(gX/J.=T0L6Q-P&L#C:IIJ.7ZR78ccQf1>,#?bV/L#cU\J5RK+P-619-WZ9
Wf\2fU.6&-<B#KG5@/Z.)AQ1=_2<\Re^SFa)P_=M@0:;>(E;_d-X785B?QR.12b(
0<AB<SdNXT18XDKWY-MCWW2BT=WU:<11&+_A_+a2bf1eX7;@Kg+8A5/87]-UM1Z)
fgY,A.0\Q>E/d/B486&CE8OJI2/?ZbWA-f:^;WM8J>IML?f+[4]RX&DF7PKPZ(W:
V:-(?G++<S^SUJR_3J?Gb#5bI1=NC>7J5DF]=CUQV(1N&YRI(:>]Yc2E(1C&5NMI
+@HO+I3?He-ZRgO@eB9+@N3f5#-W/?H_S22V>c7B;<_QKIZ-1VZ^F4#_,P>H+N]d
(64-;69)V2dB.;):6R>.3J?ICM(U/.H80\g8?>I)/]_H=/MWHUP=93HJ7V3K;Ibf
?aT[##,X:Y2?LOR9Pb#LaT1FG8+#PS\@I6/9-@Vd0,+#YKQe=N@B#>V00bJ0d,aP
@-[d1<Pd1(RM-faLWeI_QW)Ie]a(0dJ+;7DS.)&\Y;&97@X)(VQ>0H@\aBeHPdJ4
QMe0PYDFNT@A.>M;=U.,G2Qd3Q0A-AY5=K(F2,H8fc8O+._1DI][ZH:QM^N[0HQX
LT&d:IbJUg=>AGERSMd94Y7g:9EZeH:P+1N[+H&dBA#S=aWS8bCNa+gPWF,#AQfg
J3JY7TcJeUGI4Hd8OcC?0W;0;9aVXM:K3E6e;6-_K\??<G4a@_OE9d]+.H.deWKS
QU:@@=]G5UA,?3Sg8_57dYe6X&&AW>V^V_4Y^5DML#V\2\ce+7#aH:gJGSUYBYXW
^&:4HH7]C)6Y/]\fgCVIEIgE8K(c9[aYPT)Z&>MR[c-2[<I?=2-B7S)WKDNQE?1L
+E^Z#)W6)?#[=>FL]&:-VJ=N?+AfB;bPe3d.E<X#U4UBYG@L-e7-O@\YNag6+c>U
U&M2FJ<7AaTCaTA(@LHC>BW>U19U/U]GD@DCT;TX,C&fSPE8FNNJ^^TF@c\(,5&J
ZWMcfd,ZA>/WfFM6(NA@HEf.]W#99UAT2LRX)#eSCcLgcTPedFGJTN1PC06A.Afa
VMcGd)1J>=H/3K@K2@(YOa2N9.,MX@)9bK2^>f)XNC4XNHSM73=;H^T5LgfdP4__
U^#LabK+\S-ZFP:LQ&g]>T638(b)I6e]N?697AI^5;H(Zd9+f.;-cV8U-6C+>Ze<
(TVS7,B0I6^<Q40[2G[L]#E066ZOUg0HI.<Df5e/]-HJ9#M-63EgB/<(<3HL75OJ
gNQ,#Q;3.0V5-9<_8O5DFUX8\:CB[]>SSV=K:5e\7(cQf8]C\S.I&G:B>.9P+Nf^
[CD3g[XGS]:10QZ3RZf>gZ8BdeJN:2a<@J8^2G&S=0]QJJ1_D=IFcA(W(#RYPZfc
AIg1)Z;+@32G5D#I29.Lb39,H4Ug^S08CP)f_,,ZNJ49PKg@DdR^5,?8RZT:_C#_
);<<014Dc>:_4N(D=1XBa[A+:(4UTB7HO1P]=N&Hb.085>_[NMT#I@[AWSB.(J0.
99IC8Q3+_Y]2>[4L&^+e;gGd.3[#6B]VEdE(Hg(6MH-c(05YJOB[8&X[CRRg7DMY
06K=_Y5[d/BGYGU/8aJ.V5?b2BP;fK=>ff[DbN4CGLIO_.&[OWAHIB]6/JXUTXSP
8K5_,/(BQI<&S8Y9Yf494:c-91J6R(Gd3/<7R>3+B6A]LCIc,d-FU:EZX2_EDXG=
eXDPUHA;K4HRQFPWK@6e/8<L[_B+(.STI?eALI/OI/.E7,J34Iaef1DbODT?A_+]
WY\>#)KSGR]Lb54AJadCM-BaCLe&B--\?H6^+_42CD75e49&?3cJCJF7I#.DXGA9
8+48FafRWW<YG26\-13ORD0Rb))W&PE5@NLEJSB-F7RCD)aDX9/55RE(GK3]F><-
PG,J[@Y/Ea_5:Ye3UEBZ7-OY<L6ZS\<A(W@c\H\[=f=7,SaW?+]_CEURf-U@I>2)
UZB9c,DR&7[3XJOBSAW&S\c>gWHRa?&@QL4L32eF4OW/2PQ7gFaO1e>g/U4ROCOF
;80aGa^,-,QP;O3Rd/Y:4JgF59BN]0?daO3[[W<1a_2cEQ^>;(773)/7ZK4T))3Q
M=:E1I:1[17R39&Od_0BQ,eL[V3_1G&CXU\1\,OYG:(SZ/6_eb]+P36?V+D0,I6F
7HZK(C2Q]YDI?-YBb&X71>f1#&JD03)N0F,^OKB3ZgT92,S:[<N:Z3#U8IEg?Q]B
NfGX>)&M7_/H[3>fa3,-E8gA2gHE)W.MMe;_Ng+L.V4D^d1+4KIH_K\M;;FT2_Xa
ae=4&L9I62-10Q?cb3b1VC8+W-G=A4VT9SJ[WN4f]<baCS].<GXD\C:,VM1<Q8TE
B[RDNH-cgZ65bC@BfJ;d2W]=JAc<1.-8@8,+FN(\d;Db^+4EIC-K0;LB.,&(6SP8
IYVU3.@Q;RCdPMFPSIa?+c9d6fVEBW\(>]-^L2IDNf^]LUdJNP;ZD)8IDIAbGX@e
Vc/B/WX;53G0d,7TCB+(FE1@:gD#aI1P[FNc8=.Rd2I6.Y&0E^T0\aAIf/W;f3&3
YKCT;@YG7=]ce@K.SeSD=<Y/TcM5-gGc9V&eAd=2@:(HcC8./\VN&I?-HEFZHOeO
X/1U.8(e^H1-d<F:;N:<MEA9>JM])T-@J)J>7e9cQHF+aDXVZ=L];]L5E((KQd49
AMF5Y+Jd+(&+&aA5LCeb]E9QM;>_HYG<UgR_3d/00f].7KeK-B&Y,(>+ML+>#3fU
e<?E7ZHM+GE9G>f_,V7b+\1B6IYZ@MW7T-Q11I[:F_BLG\A,c]-Z:\(S@0;GJID@
V#eW5D//S_\bH<;Y]c\>&#R2a]AZAY[T:)=_5bM=^0HWN9G&(BHFI58(c;c.2XaY
)?TZFe/D5YfP]>NL3SYc(LaaONXB,QZK9O-T,A+@3_IcVZB72MTVa+/5gQ?fUKCK
_T[\ATM0Y3aXX@B3LSC3\-0J?\\<EH/>e[Zd78O\c,,+gO-1G;)I4N0C[@:a]Pe1
Y5BQ850T&?3--\9BCG)-4aQ(/gB6J>O?5G.;Ub(7<0@1f9IV[\Pc+IEJ?\B4f<Q(
:)Qaf;&a\0IL/^+\A3B:gL3&:HJTgAT?&Q00B^0TDS=G-@-4-BFLXWD?WYN).0\)
WUGb;Z0XY,e-Va.I)4/XD4]C]Q;S-,TQZ9\2I0[VAT5O[.=NZ##cHW[RS+[T681M
.X/_8?57\gb2+bU;IJYUZ7Ua_g#\a]71a43U_1Y/e)EF2[)[gB\FR,<Y91[2&S?2
F]&ZN3QL]/\.5\;,>7EMFL0GJf>W^gDV?g>ZR;.QFag:RK0?;<?K12@VS6eHG8O7
K9JR=g_G;Ng<KLQ)SUQG=XYCWa.AZAI5@C95dL8(V:N8bF>^#@D/^7N(5Vg?-[2]
5<.1Q=f\Z3RLc<XIb#6W6EGSb7f8#?U8<6ZDUY(aJJGCV?A2>>YfeEWZ?L40/;WY
.-b<H^\XH)OcJGMH\=XUc:LI\Q-.E.L-;LFK_e[956FPR+3S)T6[_;F+CD8OP#ZB
D513HC@^_4/[]JQ14CO5aKA<2f9\5W5e:N\-=70U<MJSO.Z61BFD:)FKAN.YEKX4
D5=(C,]#Y=&U.ga&cAcA#DND&4dMH7NU/7<,B,0)C-:?^,Z0XLN<b@J<-AT=M@^)
H7GGOLCR<cZL2^_J_.fFa(.:18+a_MeGQBXd&=YcSg#>ZYf5eS>\K15VXZ:V457:
./<UG<IgQ0]V9.,FJa:;b-4/A6dIH(LN^U[@HF8B)][Ba4#SLFG?gNC33V-ZX.V=
bdf<+_cS3TL\#DDZe07E8(L+d\TKdaX=)bc6Q.H]7,CZY=ZJ^]7I+KS;]H7/RPTR
^WHYf-XR4QR]g>2=Sf4Y)Ob@>>+5)5dT0EFbIXdE.V?e-;Z\#,<Z[9+Gb)A5@4c?
NC]S7Y,Da-Z6;e2>]T?495QQL&_[.KH)KRgNEY=[NURc?aDL5ae)X[5GgJS<E(&V
+\g[-:DWc8_79KR#g0a\)&a)ACYa3Pc5TS,?X+5e<7K\c+1QU>REZC7)/;7>8d-3
L7YK)\K>IJcgJS,.\J#KP?137<D2>R4ecE0OMO5GGMAA.Ze;L@S:a\ZVHEf[?4/U
=R+VM,51OUR2.YCD#P]L_],Yf.^L&[92VIWE-OBgg]bS.N)>BU@E.a3N20R,V_UF
&g^>E>2T5Qa97Q8\DEcI;^-2>93f,FE\1-f?EX)W243DOIMFBM;FYKG,801JS0QM
LA3TZG7,gc,.;2SE[?AJE2CL8OB1/4T,L-]2XQSLC+&6>SLU]<FS>0-O4SX9I=fK
Ib>B\gdS\:,7a]SC6I]P5?5\[MF/E69OB&S<0CCD220M@(KLM0#(5T57?V6C_=dU
gfc7<\bfZ;]b&-d^Z]<P,bUDE)0[1f>345L\a/W?YB).U2g>EM-OC;F31M\JEI=K
O)L9/_]H3O44?RRa@EW471BV0;I<eb\,gQZRcN.Qe.CYeb#QL<^2eW7M7^^(4.DB
Y0YRV[W_JK;I9C;VU\-YQ8:/T(>Xb9L842+55EL/4=Ff?=[LQTF-J2N;YN;S-<B@
53@e.0=755egYM[^BSQ+#&2P+29+I<R.&6)DWa_VI5fKXbDC[?L.;WI5C_VAX:K5
(K)@8>[-TM7-B/O._A_C(e:J4g6?IW7;]_U(aR88=P]+4dB4<,R[B?&+8\-IIM8<
WTVeN\+WA=UL.::Z;9W:,-B;-.WdC?e@fBPOVR8/;E3GY>BJ7D:+]\/,+-O3e((Q
0C/c&P)JLZ31P#NW552^)@J&U5,B&#_6,JG?cN)>)aHE79P;M)O;0Q&R/_#VZKS#
.&.Rc/b</e]\-?A<D16R^[<KVQ6V4^-P_34)NQ(+40@2^0dX?257<PdbSGaaC760
Jc#BELfM;VG#W\9O3VC#\_c7.FaNe6<,5e&>YXP8d0UX9\UM?gU(<LMXR6a:O:QH
CP_)IE#DH],G&?#e1+TK]cWRC[?d,7:BOO<(>=(ED-9e@8Q&T)0Mdd7IM6Nc/]O_
YD^Md+AGg@SO_8;]4\KZC/J?7XK^WVO4A0O2d3CU9[Y\ZD5,(T@BLG8;[8BQPT?Y
4G/_MYPT.I6J/,YT5<ge[AG-Q;)ED\X+cLJDK)I+GD2/Ld9?B,HYVDKG7(BX7db;
2K7PCfKL:MVc^0HFeAQ;JQ;E=TC8T&9TULb/LNI\KI3I<@V=],&/^Z=cUT-S?D8>
ORD/RgQQ,&NQ=D++<309(P/FPND:WL8X9+UPCM8,BV6PgA\a^d:(]0Q&EDN.>1IL
^=9U6b9B/3G3[N=^6Q._SG-^0,2--WVX;>b&VC_9E@4cTL]=)Te0b,N-6^R^bO1F
R:X\/1YW&#Cd0a58Z5X6Ec@JWg.VQZBP;O8:C#L]W.S28d>(928/@^#IUc3DgPVX
D0>(1+U=>LW#0W4L7(eNTDaG2/I2,ZHcMFXXc@4NdRM2dgX>Q>XCDPR-]@ZUAc.7
Z+P-eK8VQJbP&Qd3L7&RCcOOP+&/Z)O(O^=-:]VcG5SB8C3559A.2HEd3?]IC]HL
R\0N(A?P?>HX-^X@=4Q8QC[BP7#]TEZJ:15->4b.2LBA>]]ZgDOR<Y0>&e#_M#K,
7S,ZXRZH&>SK3a_3;2MO7N2B+[IA,+@dF5BT0dP2GS@2g8E(RdeP;aIGK6VgF_SW
NIb9?[]D;)7N^)=WfRE9ZJNd1]9a46:/SY8B?Y2#J-RS9AG50N@Z)5I]E/7^_<3M
JYIO]B)#>[5)RMYUS3deQKC=,Kd]#(De\;=\[R.Q=S[)1FSL3F#L+H9XF/2a=/gJ
707T<3]MPB.>?@+GN(X[(3QXG?4\,fH>??F=9=FZf8?.)E&-,S>aB2_9UgBL/=U&
2,fDTO7=:-cT)1=+@a<5+VeO=.>8;Y9S<+9R\C#JfRWdX)c)XT-?Ge9=Zf[4I55L
Y)Ydc;;(H>L]VB.617gR.Qa4Q?Z8>7fF(J1dS1@@eP&;EfX\0E\J:V]:+cWV9EF[
Sc#RG6V=E9)cG^K;H,Ad;7-C@^/&dgTN[3GUGIaT3T184X.LK\<.8g)]aKN)TH1?
N=X\[&g7L?EK33.J.8]6+)RXAF5^dY01cWc?.,6P<RI._eYZO)[^bCc&.VN[J=01
#H\&X6QH,\C@?X<G<QF5^7@A5KVf=?Fe;JHEbOPe)Sb(FM&/YP9UP/7_/>\R^(0[
/B(V&ND:.>_.0@-C]K&FcYUaJMfYZX[0K\9WR8c&3[Z20[DCfUCVIR&06a=;.5@-
-Q<TLg-(Y;GW(K6RE9KaZ]B+JJLICDV73F)N0,?,#^&GJI<+V37X-G\;6bWS@ZRR
I(>.M0VWR@<Y>CG6S>YM^]SF55Z_C;^BTP[B4_Gd/744V^])CH7V4)MXAMdbc?;1
9+;H,MYY5]AWG\BaC3_Zb;AXK@b=KRLd/C>L?HL6dO/Y7&9CRY0&^X\>f94DK0Fd
U>;dAE\IbJgY[GNgO8f>f?B0[@V1EJP5fKNX3&EfLN2O7g^(VE#CO)VW.\IJ/W+2
A/b/]YPIBOHJ^d8Y3V]gGBcPe\T3#Q4c_[#=0X^9eL26Xg-?YGc6K=A.>LP6Wcb,
5X<eQ-2D^fa[I4Z51S2E&D4d3(X1Z9C+HDP1M?aVW-<A.VFQ-UL+I9I;9#9;bF\X
)4UMgP>O./9+>d[P(D7^IK)I[IZBCWd4L>SCF)@<+66a#/aVPcG5O664F+]7WT9>
Ac)M]3>QJ,BWTaYT4@,_>R(@\,;BMTMbC^,TE\4Cd/0Y0ZC#;7/B,Pe?e7a_->2.
7J0AcWS.-RBH#\\U>,1@F.U<cFP1CZ@fG+Q4I@NX4QP&b3RQf8e;]>&_=6\PeXVb
)J9R\AgC&aU#;fRb)&K75X^BU/6-4N.ZX&6cU)BH_J;PWYXXS-LaS5AX2f9X6I-\
VZ^;EXQ+MG^?E04>Od5P9<]Gg^b/TZ-L(/L;6D^Q>cJ,[.&G4&13WbU)9TGDI,BM
\AD+g2/UBE^ee<;NY7)?H?52ARAZ?EIXa#a(XeYB9JO9ZLT8.YG6Z:BOeCJRb?X2
S-V-&dP7ICO?H5I4GEB(X-T:?5/E@ZTDO<#d=NPFP9Z=AbV&C/AIDRg7CC-8<^@]
00;8;\?bcEd0\JN6]/Tcg6b<g\W.#_6_S@C2&fW(3H@4M3IG8WD#6KNgAgT1P3b_
C,@2U?#XgSbEf7O?V3aS?V]QUOb<W5NF<\b)VCQS3e6^J6B_O95BQ;fO2aE_7L>c
+0@(@_GFCcMMU5I5(37_JOQCV)B=AENL+e5PML;DZ#ZCJZ)g49<([b\cN9\75^4S
WaA<f;9B.^?/9X414A\\g(YQ5E)d81GbW.,_;UF_ZO8CecUfNBZKL3#^@B[QaPQ/
6XP1;JOS;)QY]2]>BCY,L^[YaS&>QN.4E3C0\MH.2L6S:+#U(BO?V-5OKLC(S>Da
@/>K9J<FV7\OH=[+f1Y2TF]6bdH_-FT_c\RPeF5/RS:4U]c+PQAN@92#A]23DZ^W
[\b#dP?;-HXL@[KPCIYF4L/TTMY_JC(GLLB5OAcF90Z2@)YN>P;_<[OB/a_]aQ81
&T>c^7LfV)CAFGdacA<+XZG+T+;abW#@A>&L7+SDe>07[EL=UZJMB/AV)1T=\gZ/
<d2Q]=b2Q4e]d4<_Z=P+BAa@-NB@DX-89]LX7N^Ae:DU#J7C/XE,Hf8Ld3/4eI.Q
H972c?;[]eQK]eK>#d2;4]J_)KN[CT]VZV</8RJ9RF+2,?2C=Of.Zf^Q/)9>9];P
-KU6<OZ_VTb2e9?,^^DIXP^+[6IcA2]<T<0EQ#Ff+#OV\.YGF[aZ&)7d6d3cEF6J
75=0La&PY1M6P^0MOO;f7[Sc<(F=cP7;#YS\c[5W>,8DH>I=5KJ##/HC+ceKLMS2
=DgNaIX05T+1bgV&F_<W3J)7JXXF>>?f-.Mf#A3VZ^0WA]N;W/1N2UA#XX#>\D&V
1=-;FcUSbeCB4Q]BZQKI;@T.G;e,R(]7-D)ZPO>+[VL:SU#>WbQ6#2D>Kc/IfSKI
CP(ZGbD2J5O8Gf:GF)UO8(0M57^LG,-[f^b2X30OX8T+.WJ(f,4B<1Zd?D\C:L8N
NaPAZCd/C@b(b,5.T9_d-eP1]YX=I4DeT#.3M1A8Qe1L+d#9bS3dgP:D0)L9W@T2
_#OJ\\:KHJKWIVN-/P^1,.W+d#^UJ>G@CgEWHab_AG\_?]4NWQLb]5]g4BPa=0;Z
S)&&3HW)\<f(\FX_RQPaXO/&J<,fH]a)>,Y2&ZOMV2T\5N6a0QW3.d.^ce25X[P[
4C^#@A&faK[2^36.:PKa@/2d&LW2daE\GXU5;fF.3)]@QgWa+AE;D>CfI3E[<R9/
U\47fIDfae_CJZ?9L2TZQ(Scg-3C;(X<c;&_:(W,ggK+MN^T[c3OPZBaL=1QT6,7
):?IQ\,?HE_a^4UC<^Q\=SGMAZEc40UVeK_=SYQ??VZ.,a71N3G06\+[L4CCVH)I
58J5dK@=&<;a)<D:3IfL\4))O[QNLF72NLU/#Tf<<<EV3ULY<CSQ^I7KOR]U:gXQ
1U+#89KYeARCPc:\X?6&^^E^]Kb8>&f@\N/[+)-#K:9&O(H-GH4STea5[T8#X&]g
NdD4dZN)F?HK^fG3:fNA4U+=+>3-)IS?4c.<#THB7+??cUcHSI<8<]d?[g/+[3]^
CLI],ZN,P6U<=?B1/N5350Gd@2IAd5eBcB]<OfgF)&R)Wd3UXU[M\ggJdf-)#a4(
ed6F780dD\5T]X4?OQ8a6R)),Y83/cO+PVPf-DPR8VeZ\/:2<8#I:VK&4,9;Fc4d
=Q2./bD72N5CS@Y)A=#\KXDba4B3HOCNEURL/\b5O:>87THa93cQ/8QIRE;E5:0Z
.ZXbQZVH5+YM4ba-Q;.0<H/gGW9WY^[fXf<-G\Jd,2M0,fCMV>4UQ[T88&?EAdH6
=X]\Z_?fb3@;JW/2Y:#8)9B.X\c<5MF]RAW+^+6_WC1;4d/P:;7PF7K[T)H;d0a)
:W.PGQ\=GL&dPSfGSJ#V\ID6+_ABgEDL=9dc5e1ZZ+]A6_T[(M^ZL7L2a,?^aA]=
,^?O\Y>=b((=Fg4/^3@P]>d>Z#63)-K9ZFI&f/4H9A&1,:e7<0Y\:.Z_d)X-JNKR
RbY]7725>cRN05IR7J9:K^BPY2#W]bg??9>6KfW^V?eF+TEV9M(Gc9ESW(1d,HO>
c#af1G_#I_P\5&GeG7]?T[TbJ&dNHNcIb7M36U/U-9\AQ3A?DJK+@@1;Y0+UB)XH
gGS20-BY)P[HPJDIT+_+FD5g7,gG-_MA7<c,82?QB<]MNgDK9a.;5a?F#BbQRG5O
Z9fN#-Z,[K1D\]77D)[:O_+1R=ZOS>Z?4Tg/7S7-1GJ+Ye]c>>;>1H2-+M1,(g-d
_XLd:b:[<M@8;U1FKMaQ16)[J4?UJQY,6?e6_Jc5<X70+6;2L4-T(-8H>&,Sd@eD
>_9:4_1@4UB,[>#[b79)KI[.EYX(;C/=0N_0,U;9H@8/LeF49B7b02BX?6G2SEN9
7Y_bF0D\L5g=NLT[2IGd2Q9).Ec0;\(e?\[.Q8-/e.[eM1KdQ/D8;>[D:::583a-
BZ=7YV;&fE(1J?#,[(1H0RR<[6#]1M4_4>NH3MHMBT5#MI-ZL,@=VCN0KY:LCQN:
=+-S0I14<C?bG@J3?&QUX+Q?:,PJ,E?DD9H\Q+L6eC9;[gS>JaZFDQ4WPSL/J@[R
XI_Y_>@KDS8a8Z2aDW-W#R\_-8;Q^Rga0#,-KUfFE#c#b/eOCCEK@&(=9Ya=\#(5
6c/ecZ6DdeH=2O#U.>W4N5dWZ5?WHQ09#,7(-O[,R02KPV^O599@L,0P(2)eH#D<
NRbd.@C:Z9;11gfDQIggcYSYR;W<M63L-OGGI=-.0,P=-SBSE>AUPQ(660XDU[Ye
J[dQ&OLIL\TKHN@HaY;G,@2#[Me[F_-GabFa#A#cMU\dD\aeQ91:H\43O+7SD.>9
2(\1QM(>\3N+XgQ3FaXM8eE;?Vc1efE+5^TDKFe=N@e);DcA222J+SJ=bD+]b-UN
K]T3+Qb\]_9VRX8J8YeYK8GdYLHGKE0+BSC_^7._TPf#-?K\V^(5d2eS@4I]NH^V
-DNPeFBDc8HVHF+2fS4A-]e[T&&=U?@\<PJ:6;,VL4QXI\\[-AM^Qa;:@f723Z(6
V=<dPC20(=+d,JHXBUfc3EF#:@NV2JZ=6D>,#fLXOLZY9-Jf[&XY\0,Ia_=(-@:#
CH<&2\0MY)gS]#A#fJVO]<aWVaWA;/;fYeU#ag+P^6^&,X]4]QE<9&fAZY-eZ@PT
M+QI<0aFUcbNP5)Yge&<.&@<:>M_<8]gW60A?^\\.+.:aOfb=c8&c_ef\HQQD#DU
Ue7MO;_#^AAYce+aKc_(QJcYc:?V63/0E]-:]^KJS_?=5+>&3e^5SfbEIG+A3GD2
HE/NZR8?Xa?WE=\-N6)@3Gb2K;gM)APgL@:ML?=g#1>?+NT@D7^gIJ2)7eIeV?AR
=43FAZ;?d>YIT&E[68)YZ.-f[T[<\SF?:/1FNOE805KNdI-GYY.-G=[^Y@.FWW=c
Q(g]GG(5IU23)GNWK0F7](7CMPe&aE38X.J,=4[->01I7)LQ5UEdY+>g2&(d9c9-
O(.@DLQMLMXe78K-CYYaWfU(M1OKA603Jc@<@0C^AA-/=SD[V46]M(c+36(7L8)H
GPU5.6.4.-KK?]0N7.P3@(/W>(].(Y)MLX7HOTId66E(Q6.c@GbP>e+7MXA_EILY
TN^4[9YfWQ;DT)U^GF06B#[,eGBL\L.:SK]SXREC1Y=LKQKB?,P><S2RA>=7EPeS
b@KJd-MFKEH\S3eF:AYN7<Nfg?YTPXCZN@E6-MFcVRO>&6-@14ZgCNW_<R#&c?LZ
0:S(8:9,B,DI_,F:M071/(GYV)[>[OgRS.&S/AUbU3PVA_WI#Y50J(,>-Z(a^fMQ
8ZBE5\1OSeGK1#H<EM/?.:T8ET]eY&F,65I]Jb8TYCeb#42##MBMG0g1OaI[M9=#
VJT/:^&:3D_H2a\R#(C2,KT-a5De?/MZ5W#>8=H7F91U=2^NLW/F@CS-_2_gSR#3
a3JN(G1X\JQf=C;ecW;O5aW.>1AcO-B559;0O?9V&5;_a8^IgL6NMaKAI<;&O5XF
bSMKf.TY\&?D.QIfLLU]f&B:C\&_\QF]J&[?EN7B2^(&YcV:]XL#c3AcTTT#3g:O
LC.45FV+=ZAJ^bC]+6<U+#ZYN@fQcR3^L?P;4_Qd0F4A-5SC.AECPe+WC:TJ^&,7
e&g:G(9S_67P+Q>Fda<.?:UDP.5_c,;GJgAW,;VRU\9g:&26P-,Xf_J=Gb;b0OWS
ED3X6>VV1FC3#^8RHM#/1CTFN3Vfg<7+0\>A@.R>c9Y0Q^8H3NH1UN2C>Q]d^24\
TbU_R5gE],cQ1=>23W)9dK#ff[1,:U/W]d[DD,Ha?Z,&T7?GPM]HYA2&29=1&7U-
1=EW.Xc6IF>]d?DBN0fA<fbLMe.?>,0&Q(]]#bfc:_\[U=I@A172ZW];A0b-gE-U
B&8/L_RV[A=>IWR3eJ;-^/gM4a.WR;.VQ9;#[Z@M+QGJaYPM.]\F=eNXYg;M.5gf
^XI.(W>fC85BcW(@MfFR@0GOQ/\Q+2#3?90LXKIJ,R(PMc0=0g&#?YUKS8#bc^8A
N6=.R-YR;[.7/Q;^I2/#7g90U<TV<?acc7W2\5P,_\K^7BeE3\:c)OJ;>(f9D\QR
XBNA:,E8aB06)2F)N@@DN2)4I?O;<b(]ab9M1QF?#\=c1PV/LO9Z>Qe5bYQg0W#A
,IW,X9@].FUMU7Cc:E8JJKFKTXT.OT21AAfNZ\JAS)VDd9:U>Q5)W8-#8,TD:9e)
1#8-cgC_65;AO,dBe;-c6eWS:?8B#ddP1cRC;YaK<dLb;_C\MP0fXcJ>GW&?G;(6
^F[&O.Q:;TRW;7D364R1\4-[:A&+cU/-A^SY(GY#@=[[PC];EP7C=)SagB>\&Og?
bV/B&BJWN@VML9+\W/\@7^dR]GP55,]6_d9\6c)D#d?W7S\,&J89^3gFKfQ+RRIC
#YR49V&+V&aTXQZGE\_,[gB:;QG<S^ff(FTH2H^<,abO4Ag?P7T,8/:c:d(,Pd>+
H[Z<5Q<gE(47:_Ee;@Fe[K>JO1d[,_DQ045B2cYE-WF7_HCLaFMRACY9-5Cg19aZ
d&gH-UB+39U1DHG5Re_BW/\-AWgNY=#H>IF;;>YEQK>B:JY.Q].4)Z;=RMZb9=ZW
\_>(^F=Z(Y/>\E:CGD[fCE<g)VTW/^f.FgE7fG6<:U)bL:YSIIPAD+EKX+H4KKWM
AK.DVN@ccg+DX?eLgB[g)O<:N8;NJd@8ZX<^F\X>76Q3>.V6\ORLHFO5J7BB,?H>
L-B1dL>e@:&eUTb5J>]^A_O#XMY5<-<d?1(E=f>-_CEYb-6O9<>Cag;CYDc4G_bc
Q#Ed+aQS\e)6S,S0;cQ)PIWZ\/HUcDgUGcY<[##&IXI.<.2,7\JKIS=<QM4+]@2-
bO:S)PNJ7]f=SXENOe#N8:-f;/[0V;fOf#]D)U&W<W7[L,3fL;9APcM>?LPG5Oga
B3S/P=N/c<F<=WB1,fEK2\VVI06NZgVS<1gC4^db,O=?07_f0(IcXa+9>H_H1c0]
3[)gJ-XOR(aFddO@CE\I_S+=[7FWf.]VG^H]4O]17/P+^IVNWE0Qg#88-]_SJGWY
RE/S[X0A/R8d&6G3ZDCE0D_2AOY?dE/Pc[^QM_,3<5cAg5P&V#S8O\Z[/c(5A]E<
_Hb(+P94A3R;2+:5-YK#3QT28O^@O_1HJCVK^MVB4:G5gS_;[;K(XH+)?1C.E+A7
dD(B&^^bJ)eH[:=B]\0EM/R&HD36DC),1.<05MD\--]S,fQ99]fS0U+^(36N^NM)
9OBFb_Ke&46<?55L0JFD].B,aZ5/bZM<U#)TfL#a5]<f=^e1:@IdNN^fe6Z&Q]I4
Q>>3B52,KV@[>TgZ5ST(QD8H;J7#JYYd3I_T2dH>c]8IZXB5D:<\VFVcc?606L?<
YC_Gdd?ScC.8FL8M(dK+R02&<.PcFWaRG&))[QGfLM-7RUS9K,8KM9Z4e3\X+DPV
f2G-a>.;.?IP;PaH=L^6+g-\^6b_LZ=4&8^f@Uaa\:R0P9/c&=Y<@_TM]ce>dYS]
XI<W^I5:<ZWC.HT.&bgN3DOR:JRYJf[07LW,?IYeG)a&AE5J/_XK2V,,2Sf(T1X^
L5JZ>SQ1U1c.@&6g@bBYE^(2eO[BM:RQ?EED[.X;<NU\&XB4BK1C?57UJ2a#R1R#
g3^^>g]Ed4UUC>SgPSTPREQX3d;S]d?/&,E1^ES#BC=0-Kd,W=;4-UQ)1ZDZ/;Zb
Qe0,:0I:)L<FS<-9AY8L,g2^U&<gO>R(;7](BM/P[W(aO7])@NLA/8dJPH\BG3^(
/49;bR.6C8[#7@OE2]^(;+/+?D+5D2U?6H[>V8a8L;c=IMTW)BT/7LR8Q.6dg\@4
0,X0U>/egG8[.+[P>8U9\V36OZ>,QXL:H.80GQS@2TKBBCaIbWIG?c-+bU^+5BM6
X9d-_K[B@U2,eGR\(\+:<:[B89_>a2Ve+-f1X&D><:T^^dTVbWAZ&O_W^5HdTK<.
_TV1gTR(ga^#4,[c8PC/c+]4=@>N9)P=d9XL58@<e2YfZ+7\e6L/<eQEf=J^ER5F
9FDFY_?.-POFd\[USF\\HREN(),HC8d>AC&._/3dB;#^eQbIN4VfS([/)=9ec(Qf
8eNe\d(]G2+P\U3[).GT[055,.44(Te7c>F@]L0S?S[^G5AF>UXE=KM[]X4AS1@_
GDHQAH_,KS5BYS<Ad6^e-YZgVH9YS&&fCaKZ2dVac2P,I:D6LQZ:=eII?De_#(C3
AZ?O][=US^U(F.J?8U659Q_;PRBLZ-fLY.W,:;OG>?8#KN)4MHCC9T1B)03@K>#F
8D]U/a[bOWH=UYIZCW,G4/_Ygc@3,?RK5a]MC5APX/)]5.]B;NE#1OH)<4/=KIY7
RIN&\cS>MGAFS.U37K9U9SQP1TgD9)J&&M5_4@7:N:=2T<7Hf4.;@@T1I.M(,WOO
RCDSA_/d=IA-H.K^DS&TKP]B6RW;Z9,3J:R4<fUA4DXD1:Ecc],.\3IYMa]NR0UA
@=Z:<260U7#<H?6\RTT?20@DN0H]C/4GKcMaYQ610=eJU=T^L68\Yb_.V[2R.9^N
[#=VcfXJeFN<b3I.:,LQ@Va+,9.8K4FDN<2VPbUZ@^CU,dG)I3dg?LRg=L02.L70
_;:6Tf]DESgLe=/ed,ePT4S/IgD40HQG9I^Bg6L&A21RRTN(N.&de:,\;/,dc)M6
-:&]R=fIce+4Q6eW)<8I(BH^9=]ASg]C8JgHD[NBMc,\Z9<SHdC[aN<Q88Q>f^eU
\XZG,3.\d<G4@29I70>1GU(U935O&LKc0PT:7Q/d<K9C[afTW()/PVUE739R2[9-
e=Q3TVI.,+,?c4@EQ@#fW,JKBU]UWMQa@J33,=5La?TFK/9CNYX&\XH7D2(E.O;;
V49>_6U_geE=<YXD^/+QJI]bZ#1EbZ=Id5[^b<=U.9;cB)WQ^WZOV-9#=1D<M@XE
fcf)60P-Zd[,ZVDdafVH+5AD>X&+/_.=2.,)&b>d1WfZVBW<I_\54@[C;-F6?5ZP
3D46\2CLfJ(^-\;0\EJeD^@7_OONG2M.aV\27^)\Oc5L7#;Wc(2fMe7RVPRX\R[)
)d5&U0A=\8<Z:9fK^5BSJO3TVaDUT@Z=/B1.5_EVgL)?;:Lg9A3SNF0@QTMTK@&b
GgXeF0=X?Q8>DETKQT2.G;4R)82VS>M#YA(\ZN]:>1\#Td]:7dZbH@cSOB^5F2<_
Od+,EMF]>O6X7C.71e^PZa]=0d3M>)V>0/F:>UH^RU-+_gK5R7^c+>2>\QN]B2cW
cH05cL_P<c>3=S\O8#^@C>:P^g=B)D:QD@c2W\PY]R1Z7S0#f#Za?IZU/Pf+gY2U
dK_)0Gca8161IeQf5O7(-AC&cf;cg9)=ETDe,Yd(7a_V9-MAFZecAJHU<J8d:)Sb
SP&RVg0Ya<>_M]<?ICH4?,;:P.O(5Z;#@IU;M)[XMfaPC79XXA:@V;2HJP8g=OWH
7<ZJKSGG@GX2Q[@O3V2GYD(fQ;.O54.CW#Q<)N&ESER<NXKO&T.g[#V:f\a7a\gF
VG<g(U=[H&7U<\aZ4&R[,Jf2+,3(afIS7/D1KYId/3:A0]/[[.a^5:6L/e-ZZYZa
7E<:eOI[47[HB-T-S#.@BbHZ/J>@#)U6PO8]Md<=8O^bIZ]NdY1d@PCQ\_S4d;ec
.7+a>2_B&-UC7Cf8/5Sd+81UY6F[9ZM#fQea54/E@9[Uf>1GV8GYJ6deXe-)J)PW
&K>ZJ:2S/\UXV?C2F@/d,0P6e?W=3&8NDfG5SKB:L?7<+e6:0??dRAMc)>K20N3=
V^;UaggIcOFVeC\&402OcMDCM@-F#@Tg;@bU_Ra-KTcD+0C9PB+)V79gOdE]aSV5
:=J?D;R?MV6GW20O;1/Ja(I.e@P=d]AUG6(W#;+G?[\[J;B36X&))C,e7SeCg,O=
^RUXBf0#CN8fRPA+PW--G,\YJ]&82W:[9_g=YZ#,[0aDS09RZV&;KA/&^=@G[WW=
+5(+7Ue:QQPBCZ9IE6^)@NQFdK=4/CQ(0&;fF(Z-_EOd-L59I,;f5\7#=7<XAbSe
P:BNDH@#^aXcF-+9(K:QJ.DZ9=;WGH5SC5J:ALKASg<\OS6)_C(&P-<bL9Z]/^Bg
RYN>IX/B\?Zc7_HV&Z;]<FLe.gY#A+g=5/<7;/6;D5>^^94Y9TYgY-Z/VeIWA\PY
cYJ)F:[eR09J)&CJa6g,eV^_)RYW_#Wg30Zb,:d0K2PF2NeBC(YH;+^a8:XFL.^P
e.^#Ig24<24ZNdL/de?)>@E6a<TT>3L4YKTZS4W573<Lba,47L)<Xgd)OW]]?N^)
^FUY:NB]\)6E4b[gIYM0dS#3@[/\SL7_-A)_ea^,@GR#XdVZ(7M+a[c.Y;67EJeU
dZG[US0>ed_6C^O[XP0&^>+T>BfM_<gX,WD6d<V#8)KYVG&g]9gc4IQ+<S94W9;K
B=^]()K9L@.VY3T/c2X?VOFS;1MH.VL5S0SM5;VP5\Xf5@E0aMN@IA6,eNF<.GG6
4:6=EV<V0&P_EB@U@FI&FaOW;>OgDE]0]G[,6UZG==I3D+Qg>/YJ[-^WNI;6MdO6
Y(f\OVR1O/=gDEXQM\R&:33+R6.=d<fO]VP7NR7S#@-W@)^:.0FVB.S>[4=-f+/+
QL6d6#K)O>SGUCa1+)\F-G33FOIC7+\59U-B@/XW6>4.#FAWS98b&A10D@?b@GJG
V:D8M31T19^3g(c=^8)=U:[37/3eNIQ;29]4P7IGVY@3&LXfY\6ZV0O]5A:b5^,H
FWY_U-1(\XNK15_./eB8D0Y]G9)?G#--TMd0(B:JE)<Ba@7.(I9QVaW_HT43>>5&
c:^2FK)Q.T[KJMMg.=b6]N2d2d5/H>5;@_g1/(^#KNWUg]^R1\:<DI5;cSf?O7KN
[DI]V,?<;8e\[K?fHN0dESE_4dN-4VPGH4CgS],\4GK]Q6M[\1.:8f.EW=F)#YO0
M[OC,ID^,NKd6B(g6(@L4DIR9Fda24#dI/B0N.#J^0&bcf\5.E;HB+E2LJ5J1:.P
ObLEJc;9S]9]J4?F9\Q+>d76?fCb5-TY&:Q.7&g(FNeN:fE6F4WD9,#9O8OO&W92
Q86,d#DdL.+>CO:eE,&)^^^_d=N(/[2TR0;XO<Z+W&dXCS[+4T;:8>+FeeOE3cV7
,4]6[S@WYYCYc#RT.fbaH)==#&.;WFJaRE9CLN>H)BaA>EQB6M&JeG<IYaa7/T=(
)Y#\/c8-2NLMcgSf;=gL:[=N5dg0f0I)PT1D0I_2(L\H?UBg@@Q\,89;aFbee+&A
P:a7A;1R;Q&4WJHDS&,MPYGFGf^.bg[M[WSaE8)5P)1)E)5J@2L4d>3P=X<:\:6a
ELRAXBS[6.>7P7569S?KcbU2W6LFD??dFLdO;H)_VE9YQ<^7T-,]LQLbLQN,Ja.V
deV>Pae=)I9+dPVLH3aM\I-Te5&c4.ZM<f>R5TRBO5SB.Rc<,6gWQMFeN&FJIc:9
?O;+HDA3OKOYRd/?\OBSKYAXB6U996-6,)1NB_X)bT69\SJDZ3+-P1L<YVMSRF;V
MTE^NY<O-AAeLAUM,YNg,,KJQT5_EVO27R\gM=7V;BS/>Y.QCE\:53?J<XJ:P]W-
-DUgDbUFgb016\KHR)M+Md.e3MUF-9(VG:N2A++Q:[;J;N7FKHJ:VXI3#\)O,<46
8<F+QBYL\BK6#I\_Z\dPZ13B)\E#)YN<#8g>f&c/@F,@d5FKKJC^/6:W]c;XE/\+
;M@T(EPbV;W,^CP)d>JUcNA=[3J:L9;6B^<=L/B1IFNMVZd:V-/C8d(PX,+/6\_c
@(?U4_\-OZT:Z=2[G9ZP,ITAF=BIX4HRSKE?HTUcS(U9SK1OV?,[[Vc6O__fAXTA
0.AI\-TcU38cdK:9Ba:/8SZ1+U4WG241PHMWW[4-8N#^Ce768,EcTM2(8/S8:fcY
AcQGJ8S>0UV:858/7@@6A3SeF9/6UO_0()a8]A,HD(T5Qd4dEgX_I40c4O0;ES4M
TOBLJ9cKVa/;UfJFI66<JS;#3^63X?5-f/Y#VMFW,a,NL)=.JY2K<gK.X<MJdVP5
,R2TdK0LAf(T5gL8VKa8VffXQNf?;VR44CO=,-M>0AH=Q@Me98Q<<MWe>_T^a3U?
88W=^DX&AbN&IQ.:C7,5?IN:,A[-2a;#&NOJ#<Z67IK\EbDCD?]_KTMT:0=PPQW-
T,&T_GDW]-fcD_.X-V@^_L(1)Z<XU(ZC^H-;WBPe<PI2QU5=17Z<:8HX];M0VKc_
?EGeE^V@>7ggDggZD8eee#.3)d2U808/M?3W5C3?f(.3IG:eL?PadFaN7gMf,])b
R0H]a+]E>)J9+]2F=B#1)-7(X#+=7f>O<#/3[#QV/?0H9e_=PX)8#e)A2cdD>R48
_5Y<-/^NI=9SFG+1We6Z9(:][5cUVB4L/2:1:3JebJANDK&]I^BUK2S:W/CN,:eG
<W5B4-=@0M8eMT1HDTMMXPe^EM\[\I(3_K-X?&I1_2/U_:5aMTS;)5#CW-+d^S<g
9.X-A.Y9G<Jda7MY7bBLDVFVg&9=7FUN4.H<(,,[PJB;9_QPCQVF9T\WY6-F^HHC
#@R,KOSU3SU)fRPKEXC)CXA5.c2S0a[_H_O0BEE[1D2I,:a?Nfg9Y[HB;MXVO>)b
_F+&LLK57RP@#(#9;^)B1Q?(UEcgU3UX.U+bESYB7KP(ZC-Nd[V@RI=DO#6/6O:4
[g#,6SEXJ3R/H]/7g^80&OT>B[;OI[LF?gOHUc_\2+CCTE@=a5+T4<<S+Z+YG?1Q
@1a2,XCSK[=V<-V@LK>MPL(5QQNI^D6b_7c95UV+fVf#:2,I]3D8E8]MB.<&Mf&-
XOg6O:2XG+H7F,^BK6P7eV@7R,^(,Rb5D;\R0FNe]a?3gf#15(I:F@gM_3e>#7;a
);4JFO,eOSR#].Ra18NXaI3AB8Nd\9=d\8F<C[bP5BA<_]Ob/AbJN^e6]3U;,YXd
???\@_2f3PFKIAWIPMGP5_/IQW9WZ-Y3Hac0MCAA?@HB[[JMRbBU9eD=K9O?VFf;
,dE0:YaC>5Pe,9Pe8.YQ^EJFUggCYQD<Lg44Y73/f5ZDeP3aZ/@c,R--AFKE);N\
ZEG56@<\G>&dMTWH1I&,T(eNB]&IB;(?bPaFY1_08,3T^:7;FfN,aSD3^:D/FE>.
DC_aR/8)XaB/H7N&JVUGY+XE=VLGV(/\6J_V/U(YEE;RK<g+U+d^I,DU:UN?]gI)
1RJ).RDQ1d\6DTb1M@QUK50K^-P@:/XNWc=VA93<,/<)Q;87470gJ5U5c@WXOg?V
a<Cd]\b56^Q[<H.&.>MCdTB<Rf#.VS5W4a>6HWRQV+A/D=Q4E@&RQc4A\=0Sb@B+
3JKUM:Q-KHJ>CI[HB,g>3dY)0;[JB#6?8,]ZI,S\C).\98&UJd3/2eZAgfT>@57K
?^1SX>F[^-#5;>LO)8==1B;:O3,,S5-S[>B<]5/d.>GSA+4R0V8f?5=ICU3K(EUb
089H-K98M+^,G\P#((LO5V1J,N-2WHHQ&5=?eB#BBQ5/3;J[LKFM)\:6DZH?UB<E
B(YWg(Z6(KD[@SgXR9]VO([>MU<B9EN8RG1Ydf&_8gcRHb59U,1HYZYV-#Z1IPA^
#H=L]-N<KGMY2]U5c8=YY\,e7R50UHR[H_ITX5O4>NYED=48GC-(0<.;2#VE&f75
P76VXZ]Q<G2ff_J=Q1D.\.VHa]Jc/EVH673:V=Zc>THZB8d83,0dHbBWW^e[0<[O
[Y^]EJMI9YW@d?4L-Z5W96Y\eE6POSTQ-28)H65a>R>,efRBED=LfGQ892>QRbE)
P/EUWWd?fg&)^4ZK<0KETAX/H/.T]KcU(T&.LMF,gaZa+F+N,?WZV;0Y+96Q.WCG
YP7?+Z6&UAPGJYJSYKIN?a;DVM7>VSTf(3=&D#X9MCQ5-cdQDN@HUV3dWN9X)SUG
XW&GN<LPS=BIf=,-)3=WZDCF3eaYWYW?_/:207_^_BE?6?H6WV[#U8#^M)0&93.,
W?I3g@G:=B0gIeTa<N>?<[B)=,W8.3(,g;c\f[[MZ\;cFHLZB]E9S:6._@[<ad=?
+K=.gBPH,/V[#1[I.=/DbHM@H2TM/B0/8d,.\/-C,>]BYMNLH,U2TR:8>)E=b?4J
=4G9>8-#dK&\6W>-VZ[_T22WY7B]FDVZ@Pg<7FgJ#:NDfGNM<OMFdf#(&?OAD5.a
RaR?B)Yb)KL:Fg6WT0f_<=@RF0Z_AHV)-;gf#;/^DGU1-3BV,Wd6V2R/4T52f,-c
\2;A0OdcL2.;[R1CP/R8(1Q?PVeT(>/d(C[3H@=(b,b?V#Ma^PJbVR<d)+WeO/:@
22&2[CVdF_THcRMdM;OI5WAaG+-02V(T^_<U7#1U[IE7CV&;=WP):99D(]Gf4bQZ
QQ\:I[e&O8bM8[W=4?d_\:1;JZR>dJ+=E<CY&S-Yg>C7[J9gXEU,\Y2[E;R>#gb=
df&OJ9)K@I[UIK78Y02g^EC&T4/8:.--2P:OUFCXL#d_U@YI?B5O>Y#6>G6YHCN#
bKV/:/c>3aEO60>+:N.62N@,48Jc(f.18+da[MeP,cJ4B<\dgT2XW-C+VPFWfSeC
<d6eQPdD7RLW#7Wd8)(b(-E.UUT+f1H^M3(M>A56(.Bg&Ib[WN,dHd;1U,]R(XJ8
EJ.#A7F(D>BGN@QLEYX6KN;OAAFC^8cdY6eI21cE.4A5BX7d2-6)I3_G;1T0FBgN
)GS7[^@aL0.A2:dFgYP64EM#U@4>PD)T4(33H#g4_=RK5?;LG,f0WZSVP)70-]PL
2bPV4?);c,HBDcK[X\PR(-<BAOEa.=VX\/YVVCP[,O=.BgLA0_cCJNP7DG?G63ZU
[U6bV7KYADQ)f8fJTIc4=gH9C:]>6[-0L8[1OSAfUQ+=N2.KAgLb,R<C8d/I,)WS
e_.>X;U>NGK2#GdMLJ?^Tg2>&\9F9DH>IXg0ABN)_^HX):g7^K@efWC#L^4gKD,b
5Be=b1HAV&Q)FfJfGPcDW5d94^XA;AX9\LP:]0K@U;:&fN1?]_GWVORA>SE]e=Hd
d-[d.a^F:NXa-XT,RYa,@e,I0:1XJO+H9>aNcKA7eMTcN/O]QTJMb72FQJO\N;U;
be/8VQ:)@?Z>U9JLPc^=FJ36;23,2.+EJ0O92OUEB7@LO0)>_WQ>SaW2MZ6G8J=_
d/.,H&gbMa(Y<29c;MdHAI;K.;V\)=#+gSaN+@L^YSMd0S:<V#YN+f[)cfeSW@V+
\W)-bW[0=fE#/e_c4J9:;cd.>/:BB?51[UNALSB/U9#OIeQ]6QXX.SSf@RKT/2U/
P#+[01I]CbOWK/?;3]_UI2;9+)KFg[XAQBQ9BJTPM-eE=N->bO1-PV+fR6Pf&gV,
7B6QNSfd)S=:T(RF2.\WR?6F-/R-bN,VG,=cETM\7HV,;Y?2SV/5ZV0eS?.:J.Pa
73<F_gBHUTIOEAKe:>[13EHBCVbe]UOEU8@X;2.7^baBFKe#ReL1,[[/_KU;=WXg
Y?NPBT9]W.2DWD:&+AMBLL,6^fXN8HG0eDA&1_X)ZGR[TWfV8&^c3[AE=XG_CM(S
)ef>()gW+_U>?(B[;?O=4^33Y=CZ(8:;-,GEa=?UR<dHDM,:6Y,1NQZ0bfeJX+)M
L;2^DSK:T9SL4U#I^+BTR@.bAdM1I+X8WKKVPeH\6)O]9S;65D]-Rf;6K0Y<3Y88
+5QU:N&(NfBdW5;]K6fRRbPR/X(@-G)S264bGf9?^M.Ig(KCR,dVBbPc_b:IeRNB
fB&#fI@>J]_,^HK]NVT=?K3:H7JgA@A&W#-b@9?=A;HcI;g(4:N?K3UCC;.BW.VY
3Q@U:g]@&gUFI-1N0<4SK:cAgB4JfB7Y+/-FY:9RTcU-#Q8+>F1;7f\F5./EA;?\
?\X;5FHZNeB6IV/:^:;C0NM#P\0>15T>R50_NJ([HUA47?X6>eaU^WL1F]]Q)Z^9
+\>.VC08?Q#-+&WEcc^5:E<M-#SIOf^e4_R6PAO7Gf4YaNM)RRTBJB)9\Og+Zf^P
?C^egY1BYQUT]]^=?#30L+^67^0W\B29M<OKLC]3<(g)H@MFg^F9V=9>8@_OXd)g
:KcFE)K6]:33]6BFCMQ1V.S(]T7-&>-_0PM&=a49\Mfa+3C95D>g.3XWW-3Rb@0J
X9V,GX>_RPG;OUU6PAVdZ^_6FR)V6YT.,&[D9=V38-K.1J4@66GH0ON5.aKD9B)J
XOEAB(dP9W86XAB4fI5I]>]HJPe2&a)M4FeNXbb7E+cbAXO@>#U1fO(>_WH&DML?
N,Z2-.4<Y74FHAdd2W,ZY&#X<eP#BE@351((,L,GUG5Q>1C[&C9:[(K23cHEd<2?
4W/TIICTC/TcIV_F.42D7CO+Ya\JfKQ6/+;G2#dSIY7.e1_5)_,8QO7-:/^X(@12
6cEDE=)?Q\0Sg;T)g)aS&YO?85D6;=]<DQ0&3W2>\4<B3TN(_3[L4N2,.I,XHGgL
J&5C]0D7SD:L:-RB41-EU>EgaILHWT3??O7ZgJ+@/<L62<HG(#f]T2?I&+Ng:P(9
/JMQb=T2<.2G-)7K3;@HbU8dY@6V]OS^H+,2G8+e(+CeVLJZf@?Vef48Z)QgV][7
FDQKVdbH^L&/RV@\\NT:O\=1YY)a,6_=IOL;RZV,&Z)):>-f5M1][5eRLD.#J5ZR
ZNT:T]4FS?5/&Z=D)I.?c)3I.CH.g=_RJF_JH3OEGd:5.@07:M8;2B&0b1<=VG+1
cYZfeD_6->YXS<&F=QGM3I\W:L@WW)_Mb[Mb>;HD^<Y.Y\OGY/fI@.-f7OM&XXE]
M<#1e5_U0YY6Z5;1^:CeM-<49BO46FK\^Y21CVYOe/S;#.V/K<f9>YdFXW>bEXgf
EPO7>Oe(\7Q[E=\H(-&9#fA>ST/0EK<Ub7,25N:VAf;IH>_aA)<#PUNQ]WR13Q07
2>;3G-IMbO6[c[c2-.M_O>3B6ST3O+8(P.-^&L<Gd+)NV1P&NC>Hd]C)T@-2:&E;
=&Kf[J)\8H7WKYb?VK@;^.19#1#/GR@_T)FO[G\PeU^OWYNWdM1e0a(W1VM_Y)DT
(1P5+1)LR20bI1KdX>aA3CDT&ZTda^dXW)8+Y\R+@Q^Jd+_Id.,4_CPRS)U^42@7
gS/09S44fNK4J4Jc083NK.UXRMT1?PPH^KD.9FSdZY)aUQe0XI)?D\IT.WU,/DHg
Cfg&I@eL9^XG@=fQ<+f=aG.S:R7;BGH6JK)(AU[868.,Z5\gA,<\X3D:M])E6E(3
16b1ag4H_WKU6f_aC<P8;eKb]#1>ZaGOe>?Db0/O#QWH@KU/2AI(5N)YY;[;ZeM7
@a(/&d4-+O?618.UME211SO99M7QBMa3>SQ#J<3Q[WTg8AaaJRA/BeV9-JB^7f:&
2>WXOSY;B?Z3CPHAF/;K#5b>@bS6DQ@1d?dJ/,A2f;M>&aHJ5_GF\1&3?>Z3ZV&3
&K<CA+D?D5XR+LcWaIJ\)HTWNbK6[0A<JB0NW=M><ZJRg<PO+::XXM=9QaSDfND/
f)CMD<:F]@KY35Z^E_BC]73>E]E_b3CeGcERV[NQA],c&X00/)[LS)7U2^.Z\E8d
;&)(2_R/P0Kc1V(:[CJZ#BE21SFR4A[@dQ5_H3MST0>D<8S^L0N^ELPX,K/WOT6d
]fSB=(7W0]-X\_ZY:2[R8+;>MbLGBfOXE+GL[N=&<SSCAMWdJRbO@A6,<a0U.H[R
PY+].R?aF/2KW^7dJNg\W8;8f1+Zg>G6H2R8?)\eHPDb,4)b)(PTW+HQW\A7[VMW
:)0SC:Q1TST-aP?^acW?Xf9@eg9397QFWSH3_d.a8?U:GB)I/S@NX,K88[Y,S?]@
W>>ANUAS_Q(+OEbdP=B.a@AQ)B@H0(U(IAa@d]-de\CV:)^II,)6L&5EXXdV,V?0
a051@_VZ.)f-IE@UUM0Ve<F>OPdgXPcgP[_eB((:^L7B[IX7#ZB6<AX12ceQU-C7
O>5U2:SO]Sg[TYX7LHe;EX1B>._0;LFM7a7&O-[L2PJZ_-M;aP?=NLY97<dGZaRc
X;P][R1?@==S?XY(bc1J.LR.C/B(0UW_CXdI@W//Y9;.@aUXN]##,+D;MLAVb>E/
SSV^2#Z(a\)Y[W:6I+?(@H7RXeW+HQ\eKbgE:d;&<-e@7^HQGH4Y4E7IOaD.<88Y
(B\F=_:b7b)eK449_>Cc=AA,HF;U:8[=We>?,\JO@#<JG=HY+N?,#=X2+/M2E8LQ
LEG@6-IY8<X,JLQ;@,@Y.RO[W/,F6<X8Q)_7_UJC0Q]..>gKO2_Fee[6[=RZ/8D+
dDY+5eZ#LXa_DDTADBPD+MG@<e@]+12b)YaU;&CK(A?.0_[M3/^KJB-/R1@N40Df
P1PMd8^UTA-7:2W42\I-BUXQ6LLPbXVWK(.T4Kgc?,C(b8[b_a;/FS8FbQ6@Rf[7
&Gd^Vc8_[FV4C?]CW1I<;CJ/VB:+aXLeN3)]ce7L)])MS@+ZST#Q55&7_8VOg-<Q
G[J4(FAK1+R]8VKcVV,JR48b]AfW:e-#c_1L^JTE@.C;GVB2UW?GY;ENRB4SK_;g
K7O\YfOCSYVGF;cRB\GSfI9K:DgS?Y<ZT7BL;O7aWU]@D]H30a1[N._&C3cQ(VOe
O5,/WM^JIG76XCPI0.Z]?-0;AgSQSD.b+8_[\c+A0fW9g]IbBG5SAX6\^fdaI)VH
2/_:9FJZ(C?WKL4M;^4<I)Fc6431\Q)K?8C)c;,9cK&..6CFG2>/Qg1^2&:F=T]B
L3NF:1/W0:JG+;=KGbZ9LO:5@6I+(^B8I9)03eB49cJ4)^FLM9VCL^ON=5W]LK+-
=:S7]7KV?/-?bI3<Q0FO#P5L:;^8I^5@;JNNE/Y>_#MKDe<fSCgd7(V^@)Bb^UHD
BT99XAM[R>D[YM7FfDQGeY1O]OGcU]MdBdP8_Ze^;9g0G#0\MY#-Af<g,;\JHI,U
(V.dc@4a^>Dd4d9^Sf16F)&S1:072@SMY5_CCCDg.YPLJAJJ,VJ2gS63g:7D8HKT
N3.T_b>#EU,.]CdO?,EJ(6MK8RT<[\b9PVf)(^PC?IQNU[[160CD\KMZX(@8FVGS
0DgUT_ZF?1Q_Ya1+\(aWS3-S<eb:S3?]/Ke[E3YR.YT6H)A&KfD1/1O:X?93C:GU
f0)E6&aL+MF-3^,<1K>L>)(5N<+9S=JDU4>Yg]:[g-f7II\_,]JUJTdP3A;[W5dS
?=a0I0LO&GY1W@0@3;beRT>)J9P]04\d?]^A(3>DY>>\GL/.NeA0,2c=EO_,2cS\
ZUY57>)I:be3TG_ZH,,?D/_JJ70W7d_I7&FP3(J=JXDOgTJ9bVBCEB^Y7];OO[3+
K]_U3c_&H;Ea3K)[\(9+3&?XI?bPa^b[+BKd6E-eBfY-c+;>38,LEB)d&O0Uge-L
M-,5.<.VFBD1T\15\L:UB;03U?SM[I9RG@c0Uf3(6KV2OMUA.MPYH?7Q[g&&(OgS
UG5]2R+W>TfafF]COc4OAg;I48+B+TATM2GLd3MHB9/1;,2AVZQ&[H_ZHF@5,cfF
\]Hc1IIFGHE.Cb+]@8#GUW3ddM_6KMBO.Sb_CgEaCeJ(>AcQ2L))bQU&K2@/Vg)d
;33S+<aJN(DF@XWC^3CZfU7NQ-80)A.(c4W(.,ZW@Tf^X,EL;>^BM3c\L?e2eOJX
/YU=M>KELGZPedJcD=U65F>&cAYDZMAKMf0HYAN&WI4R1B9HW>ATCS,6[>]XX<5/
Id_D_&?Y:2+N</V-g?-,<2/@V13OK+>;MC]b:RcDBffLRGRXUagaJ2d.=V>G@XIM
>Ocg.81egJ/\V(D+/g,6Wa^>M8?5M>I/ZA8JS)C23?MO+Z5=,UQ_ZF>RCDa_0V_V
@[#;,0U[^_:O6:\8a]B0S;c.b@g4)dWQICOOBRT4M:JO(YU,b:Vg9Y8GHV+(LLX=
<>8bZR3Cb_X1DdTK<ID-:cGN6?4&1_0]/]88SOT8&dLBL\Za+-a^6MIFTf]JM:>A
V;17,GZY,YYb:KTI)_I^+K=JK97,dJLZ4Uf8aCN9P;1ICW#Y#4W4IYc6AG;P=&^B
@a)cIOL8,eE]6W=^Pf_EY=PVO<YH<3.0KPeSCB\+R>>I\Q3_AeYG>ggFGdB=NF3?
EG=(Tb-NUQ1UeM3QB#.Y<PV^JP,Z>FK[;#e;SdZ:^fJ<OfSd&DS+d_Z7.BH]P6^F
2^e._VcdBA=+AUW9N7@2/DF/RU/PGVOOU5A3QI,7)VC.^ETcW>^UQ<dLS/?\MN\:
ZG)7:VIOL6C)8DN1cQeH?Y,,M9X3?TU230/K2LDHXS^YY\aPRGKOL_389MU3T.eY
0aMJ-UDZg>_U@(.7KPLM]:Z@S?TRH@W0Z0^#&5-0W/CFS^cC4Z>Ec+I,<-O+6cbL
BT]1b:>MDIM<.[e;-C\-M+J5eAMRU?N@LO:[J(63c;&AP0_K8<8>;7f5:?><VI0^
)\JK+WXUaN4=O8+BH5I(f^M]^4Z+CJ,:=0dJ/3^S=IGUd>40^A^P6L;g)\DgRFVT
SO:c?Y<@:@?ce3Uc&=07Of>C\OH?YC+=)JNCN,Z_S:QA.&BdYNHIOA#-[cU+F)4\
=EOA-]\QecT,>_1SGE7^H#De[]\6gaeSG/f&,84Ee-W#AB1>ac?R9D_S0<URLZ/)
4?&JBMT;RICGB7K=Q=;R7;#V2?eMSGX5W)?Q?N52De2I/@dC&CZ2fe+7Q&JJe>HM
:b#23Q?VcC8FO@[B9@1ZWE1<+)P8E^9IBc[eP\2P.gBMIY8]QV2#QN<0G3,OcCM9
VO+>_X@_Q_Ea_TU4PK85KKPdL,6E&@@;6R5(7BbW9;XH,eFY56db#Jc:__\,99>1
#5:aW(2))d/dVS5(&5XQW3F<XI7d345CNLYd)RZI?]9PK(Xe0778UN)Dea=:eGcY
;,YIZ_F=H78[-M+.-31E5bYQ+;^V?fB[X3;2Mf=e]&cIP:/B0BVBM7-](ccY=M>(
(SLL]4@V]ZR4M1NK@AGNV8P]^PaCL(/#&X#/g/\92D8Re\;fJf[b.895.\3]=:B-
c/CGU9d3^ZeQEXV94X=;V?gMB77_\=D^CCVG2=9FIVgS=d_Jg.f.I&7&#;AS?.K<
]E:f:(a=gJfMO.ATVVN]dN_PZEALU5\]TMg_c6<(92:D//OcTFH)?+FON+WEI9+?
Y,Na;_AN7,.5#X.d6N2g[H9[SIS<[S\Q#(W8;(?VFX6_Bf5.H\1^3)4A#(W,Pc4b
KN9(8K?&27(GAD=aZ:dV45OP>]=LT,_T;f(G1&>)D(O_1)F@V]875)9U)aJ#KK21
Yb6E+X88,RKK(3H@(VI1/,X8>;6d7\=EDGYGc<4IaDXdaK@>/K3UdF#A1DH(Ne28
Vf,V1WI9=F+/D263>^BXTgd;e/3:WR(Gd-V@ObVX@AbI,Q<;/f89&&H;]GEJW/OK
?N,-DDRR0U?baYb,YMFI/RZ[6dS[0a;@@<+aI;g0WVIaE=7cCU2;#O&I=>AGA._c
/G/-a7[C81ae>@52dZ;Z6RVAULPGdJ((gUgJgH=:W]HT?<C>Ha7f^YFcK;^g4EMY
1?:B6ba>UXd8a:D#>L\I0XC_35@Y[>5A-GY8]D&UQ,859fdQL.N&RW/J6?F;WSO-
EU8,T7Je,0^eM24g[^Zd]N9Og[E&P^Zfc_GMO^9KbOQS(#@eIP#EfO/VXR,FEYeU
:ZX4ge7^PUM?UBSHB9L=b5CMVW/+LNL^N]9&YfB9&,@:[BN3;U/VSERB1\I0S8-C
-)L-Tg\Q,>7[HZ?]X5Ec\fbBRLC4V?R\T3:T7TBU=2dQ#=.1U,\VAT3cgJOX+Z)>
4;J=^[2>dE(e\eGXW.O0OT\9=J9CcL@2WdEW@ce(H]=47:X(=H]>gH?Y6K\7?ccK
f?:6MWLABcN#d)b]+V->#2(.cY4.S7[>Z(3[#,V=2#7Y\bE=_FKCId91<?6/>KUL
EPfe_LRF,a(N13RR#@B1<X27Ac;,GeK6;^+<>1?8[XDRgM;EbA&#Lb^8H&d/6[@X
\H@8g&X#I?HU@FGSf0a/<MDA:(ZOI[.Kf0X?b-=U2.Ke=0ZMZQ:JdAS5#f17+L7;
&adUQNe8RV,egH(c2Y-_IcUJNB;TQU2\6C9cFcOMb5]9:])_-]&5Q4+@FOE&&S^(
Cd[O7)1gN<3KdbD,&6cf:JLE8_J3d1/&WF_Y=-Z:9OO;\&ED=IZZF(.FFM;6OD[@
F9;Q&8K(E=X]QCBf\gT\Y5_;aG31O57^LH]HL-XHQY2RaI>PM6g=Y&ZE9HT/#?0E
(Y=N;7e3U1BKL04FM:U2?DPY0F8PE.b^TNF?\?)A[]FUBb8^U?Qb13F8GJ8X>Q+0
U]\?M]2A)]^&ML>T=MSL#4ESEP3<Y&aCDC^:5eNBDde_YN9D4DGD0WWMAc3_L3=4
QA8>ONJ?dA5UJOF7W.>U&CS)I1@8&SQcdO(BFHOXd-1<ZbZJ?_6G_=a#Hg]IKV6b
03(\N?0e00/8KQMI)/=6-:<UR^D/?W3T14D,1dB//b4NGYE28396G(TTS?9Y3N?X
O98O1OPZ90PfEb/Y/#TaeX=\#ggeBLB[F+S_S_Eg?dH#GD)KB>-Gf\d&YNIUF]dN
)J9HB322CO>3O7=cV:FWW8J.I3f^YWL;4-f[0A,I2]@MZUeVF2Vf4025H[NGB7T4
_U[\FNDY0:&SKZQf+G(_7L>WI<BQOa;d).>gCZXS@FB6f2/G[#[]EMC411J+ebFV
QG;ef]DUD\b,WFET9])T2OKK#dSd<HOV.XYY+6aG98b-=_QOeA-f3:JL_9Z>[QPK
>,S&1J1)U7-&Vb(X:@#1eW?K)[_NLFH0[RXVCFL(VX_D3Fd7KgR<bLO.3,bD[g[K
aL[4X.]Q59:1QW?/Q6<b?WF(c3S.YOEdg=;,^&><->8R;USfX[>L.3SC@K36.gN/
X@cYRD#GN&FA8JN\bRaG-E.N=d7KN0G]2J^8X[2aSAA_]gONf7dYEIWLC^7HO<U&
9&R_\UMd@B#Me\ZC)/aMVAP6cbP8d8;.QO6#6A+Ab=cQWJV:5UJg4&+d;b=X@/[_
ZW2ag:U42B&[T\0;0BW4=F&[\ZCL5.3/[-4=Cc.YMP,6WP&.:.=W;/N;VBMWE:B\
3#>J?:L46.NZ2[ZYGM[/,YcE8+M0[_YgBAOVD8\)Gg(ed&7JE]b:<gG7(ZLd:1H.
;W/COTe1gcS16^0&YRSM-+G(C1-6M[cQYU94De3)R]7HfL-IW/,\fP2#76=B_(8<
FYLQPIE2X.e.?QNfW1HO<#Y)fLE>.1^)884/b&@W6O+M7XPd.EgKP4>6WQQ^7ASN
Zg2=1)]NOHIaLHA9T-gXR4.-12LdLBB4W(dT.MQF>D5>?[;U(T3SUf0+H#PDW8Ld
0bD(P;f#E_ER]ObQREVgcFPfdJfT=)LET.DPCM-;e2O.276gG(/?J/JcL7^_(gB2
3aeV^@9Ha)a[d,@_2Lg(a6+dHUd+4<KLa+Kc/YC9=O=9/7#T#dX>f>Iag]Z9?WeI
5E>Bf4>K=B0M@g)Pb6M+/6c[Z_\#/c\O=(eY@XFB01Ib=V9g-O6RQHNFGfLV7G60
VLYH.QU>/25]6PgVIC2,5@>^UdD:Gd+2;>I8DS<60F(U;9SQ4#;+<ZL,GcCgFB:d
L[YRYZB.J)F+VWQ.4IVFBZb#J8e#3RM+B2c1>=_54(6.(I^I(CQ)&/3WU]8NKX)2
>0L4Ib;/FRc-/BZ-^=W.WO=&]T+V@5^HRTC?I(ZUH7#(CFLfb:O>(SG\3]ASW5(B
@9P17818QL<a0+-S8UM-X/JN5T]GbCD4L)@7+]CV]D_]V?TL#?S\X#+BY..KP)6]
F/61bS4Z?fL+6-GN#Rd(/75X[-PA-KSEOfTZ9B)c,85E],@g\ZE?Q7;bM45S1F42
?CdEM7K(>2PFB\?D]HMD-C6LA=fDHDCV&4bXGK&J\MfU415B?>6f\LcbYT&;F(WS
5PRc=/>:/7ZT/^LVD2ZH2d,E&_Za];XdRd:JVNGa_X\_Adc?IE2W.DfI)EQ/;KY5
2>\F1?dQZB7D&SeaM/bOASEY.N][;ec1@S9a,?6/^^?)b2)5KME)O#QLW8(N6N,0
+@JPV4JRbIH3H&7X5[O^NOe()VU0X#<LcTcMa_,X6NB>95M)1CC]ED;&4#9:&T\^
3\D?1D/<JDO2TR,-R8c8,F+(YVRJ4ee)#I:X(Zb:_Vf/AEA@&OKSbP8MN;0/A52F
<)AE&X#P0Y)dBA7,1ZeEM5VSaEG?D;1#>6^1CGd\9&,-[@VQF]gA#K;#J6_O4(-#
\8g;&3Q2M)#Z8[6<([+L/VX354HG-LGTNN:54UR8]\2d1(;P?1^)a@DJ\2FEFcG:
8a7I\=4SP?/?S1&);NS7KB6RP<0Q@Z7B:Tc^?F9>)-a0U9[WPE[8cH<18fL;bAda
a/\P5\:c^b^R9^)IZM8e@YM<(;BOUQV4TNE>^[FQgA_=..\5f@LJF:P#/.HVKA&5
:)?AHc.e5Zd>^/-0c6?#68(\Q=G6><TE^Vf4b?7+<,6E.[E:HIT(f]+Q?D8:&BG-
P?Tde1C9/aa=6PQf@4FHQ6_EB6g[=Jea@E3O<9DI]&B/+C[\+1_F##35cHX>T))f
9gHT>,Fc06OR\aa7XXQ(DHc9I5/1,Pa;a.L078b^7UQE=257\B2=TNQS^,GES(KN
I>g>VHCVET@>Og>ZcY--bPYV6.7AL7LFEg<?[7B[+8L>F+6A@KHHC/2KC_2M/;\Y
T+ABJd@deN^KSCNGPWg4)[/_35P2KDLB>-X363]1G(dI-.DWAb2E>Hd]Q3RPEb0e
?c2XNcSMLg9\,FT/1_^Z50\Uf3IFM8)#,,G[d;2+\[IXSFW7JF(DF_G.NEI.]+I?
)&_@#S26d<B;^,J4UJO0d/JOAd6L@M3H<A8N;Q>Q&QSLD8\LPd]c].b(V+4=Y>Eb
Y7\2KA-=#c^:H(T/YQNLY?AC0TQX<d6DJ&5O?ZM64,Y0P7PK4QMPRZ(e9K]:JZWe
6cL,7X][N3DVJeW]ZRN,XV);7cB3b[&f3R030R,X&b/]Pa)B@b0Z\Df/++9U1YHA
J,SQ3XEdY<2YU8DE,[&dCO^eE?3Q1H=DaF/ae&EIA9DGN+0Z,1<X]2EQRa#Y5N)<
1cgY5C+4D)]&8(;2#1,@/-NM)BTPf1gCQ(RZ4JAZ64H9J]F]A@BOEOM)Y&<>DEX.
_:<Ng7cOJ+=<RK@D1SXa3e-(H5UdFf:44TccdQZ9PAfOdG;IDd\a-^Q55#B-^30<
WVHHR<G:OB6g4-5\]_\_GB/2c7G9#^UPfI4^CRO8[#U\<F?YP1674\XV2RDYEPMQ
[4301DSD(b\FT7896;KSMdIVIf\&I1Ge#\?26?#0^AQ^+#O+KN?:,;8WU+3@?VaE
6A+2-+)^.2B_//ac@9^,;?J,(BJ#)FcKU8Lf\J7,VCcf<\2V^/Vd2c+ggG.HaMN#
VDRfJg__b/OC9,>bHa;.(5a[)5)]CS4I#aBM<4BH&R-8M2V:7FQ5,<K9:ZW#HfT@
CCebLIYMc9XG>b5CY]E\aN@JOBS@Ob,:OJG+,e775PY_K/#^1RJ?/W^D?=QOK19c
_,5<YBa4aA6<-^VB6BRb)Y,YFQ#;d(AXAU)H(200;F\-G7?0FILd)R[JD-JL.WAG
?2VaYc-5gO_K&f)b\9_S6C8cL4UeI^Ab9A0L]]J8_?>6;<<Y20QEI0dI7:S7c-0A
>(.d(MD99H.]<EMTa])4cRFBK-(0&@d01d9?b3b,[9Z>BBZ4TJ:C.Q2&R&IX\:O0
JeS267aFSe-=fJ+OPCZRdZJ7.XBE=CBDbbR79fCGP?f>3L2F/[L>.Q-7H.g;K\Jc
/>AbM696HTR(10_)1\79bC&0ab#e8[M3^TVBU6F1.M.<_V_K=Ke[f1WP0VX)6c1]
[DOI+(=>eSc6X=eXZ;A:(egfb_@FZ)?]+KT6I8=59e8L8OFUS5b.NBV])d/DM.aS
J>,?)_+BNH.Wb#]cNaQMQ60IB=gV==L6G=DI.98<KS+^+59COZ4;>WW-^#GCF9MD
YHXdeDVB0:aa;bW##eTOYcLKUDd/Ab3(g-J_HfbPHS[&fMI,aG+f]E2T)aKSWY@M
cc6:6V-40f28JM_SL[QQNbPUOG[\^;;CcISS,gS:E@)R<JOJgc]:&?P?I[=MdP(G
)RD,_UL;E037.:Q+HG/TC[&42d;8MF/.>PI-KZ:aXAH/fY8]ILB49LTC2)D5#VGF
/1>QZ_T^I/Tc)8f<&NT:4#M,4QZ-YM8#YVJEf:TTHO:eJVg=9O4JIBQ>2AND-&;e
?KCO<DXeMA2?J34-S.M&g_]PHK3S_(X:A0+4TQF_B4OM@VGDCP2J?/E_01WSD6P8
HZeM9(P+[)(b76.14DYeMfcS)10GB+C2ed)-R>.=cV5\c?c&9a_7NaI-Ke34XP5F
5UF4d9#FST?Gc)6T.>2.>0SDd8L,X,G=fUNM82MRb2@]c9BbWK-b]:f4eGC5-@H-
4AJZB#0N:/>/NRf=X.\fA2RIX9.J@<YY/.f(67NF74CE(5Gf;8V)75&0e_09M59(
#cC3Jf<,DeB#U.+U41F,S0ETY6D[YUYL:gaEI5d@Y=].fb0QVU+OC1QSSLS#Q.&Y
IZc,?aT<G6dVQHRR(1LF(U3=IecTb.UK-c.eM263]QNP3#bd)9aR]KD=68MXeLF\
9;B93I0-<J>,EIIFJK0F(?VdF0O@=(KW7[M)S1&dA,Xb+^D=SB69<8G6;I>82C>L
V+);0cfXWE7LeWeAVM)@D1KGP=9OP:\T>RQ/WZbW4?#I24)LE@VX-6+ZKEe/1D2d
0XCCdTO6/FdcB&Df431X#TQ=5H-X:BO/T6dT4A8@gUe;(b7UJNS]NH.,)53W?-;2
>IHBKV,B<5WKf)8/gPEK]&>#_0=QPJa.F9EI69R?7/ZP@MKDV9@C04I]7L\.cHH_
WC_2TN/\V5T#1.E#&M32#NVO-THP/S3XOP?cfKcUV1X<O&XH3;.^<0<0\_&18/f)
2><X?Z)a6Y#@N^=+YXg8)95LP4H>#(64U&)[9d8/PVeY4Ne:0AVIPIU3c+eNB&F:
fBV2Td.[?If.2WTX&\L6;U[4>T.<KVMZ,>/K.e@PeC4Bd;G&)P)8<:^B#c1cHO;T
6\g4BY#[/&YHa1UA:fCWNB4N/N@\CA,A#WaF7+1C3:2OHI>eRc^QeU@?EQ;7BM2a
TOT(CW)3],g+?6g(VH@5aFU\DF&ae/W(YGdgRJD-X-^F>AVOHf<RY,5X(-]M1,VK
=5(+:5Vd6:=>1b#8d50<BTB8S_a2&N#SF4ZLI#E?DYaJPH;N>(Y@dce8VZXB+<bg
5?UP=bL>CR\W<AFLN].>bQSLF?YY6MEPdd@1?@+cUB77b0.P65UbOg9Re79,H>;V
&F@K\bg948.0U))8V6/Y4/J#eCfO_P.[WS&?ccI@X-e<I@\T0R4/D?[0GTV7J9<N
<X@U_BU5^A@@c;d[AEb88A@d1V?],1FQ<C5VMEdU]d^W8W@SWg<?\GAbCP.d3d3<
gd_afB,?Pa8bNGQeF@Z/W[aIR-2c0b?bJX3U222KAOU53\L\Q&^ZDSZ_6;<NO<(A
I_CQc:Q)QK]^d.ELRQ)7EEgcd4:8N]a#4)[bW3\))C4-b5Y&.#,&8(3=3dT+3GE7
C8FS:Faf2dd+_,59+=AcCKA:gAC/<-[P8=NY5R2AF5D25Z-d.^I(dH>_6MJPBUUD
cJ/?cL_3Y+WT/[63>f9_VK7-:Q4>3]#IYc&7OIX3GR[YaE09fHgNc_dg72L9ONCX
f^YM.Q78[U)[V1(_OE-:g<2LENbI[]Ige8_CU95?8U#BccfO(#^EUb5&;H&R8]W>
MKa)CB1JE\gFO.9>:</;9E.B1Z:1G-c;/7@@4)7I,=/192cc9R>;-X>;U>J?Y_)^
THQU_5/&b1gW#H?)U@HY,fa8\3P/\X26FeMg@@@(;)T7,;YWQ;Dcd1Q+CZF5I+#e
gJ#8G5b//00P/NEb2g7W,ff0)@(J_?-4fF)WPgb2Q\H_:M<TaV\9HA)50H&/eG3,
T0]ONR^aF_3LC_A?)eUBaNg?)ZfO=f5X1;^:M^IHbZE1,WGQ^fa2WA;8RT?([8g:
)KQA6Z##9FRX,d,:]?83(VJ1ge2KK.Kf]]eDSU&69YA8G3)MSOS3d-0.G@MN,.3-
D(5A3Ga_P8)ER1EI8LF97^N0E\6W/2KYK7Q,VTcFZAUUB/+[\AF<Y9U.;[g98d\Y
M?TNfKFJbA^:?\;e:QC+_5d05BF(5:C.C?eLR60>5NHYTFU3Tg/.8eY77MBR=R#X
[d)]#&eZGTT68Y9dfPbMWE;@.OJSG6CUHM9[CYR>WS&S@HId7_Q35EKg9#;FR<@8
RcPe-O#Z_a8+f8_#9Ng&K=f5-/YQXJSV:@,^85B;1/5^b[?-G-7DNEcHXa6R6XK<
PAB([gCHTM.X=0.@.JKPd\MA5(:?L[76.2d5GR+C?M4.4dT.L7DP#WD5V7=1C_P1
[9OJ>_4R,]B)FA:3_+(C4Yg/BB&SVFT]S>3VYJ\D#-.H@FI5:(N3HR,(;\bWfNY3
W3VO\Xa_3O9R3g.GF;aKF]L/QQD(0-):e.HL(Jb#aaT)22/c2-eE+g8,42Q/M&>e
7cHV3<C(A+5a-E,8_G/&+/=-N#5e5@<IKD_X_)LU^KJ.Hf1=@=+_IGeHSJY9N28E
PP9GH^6dKXST\a2gJ-^IcgRAg+SW0K>D>(9Zf<Z)<5<V(P@REH0U+9?ec6\(4\.[
/73W.#e(N3T;OW:Q6g1MLXO2bL229XKIPOJeO6c?6T5\2K>\BTeU^(6aO&P.e#&:
>A;EfaPQ=,OWS,T2G@W1I(>IT>:7b8@:GCa/2b-[HF6_TK]MA]7B<W:\.,/5C/BI
e&f6R1UZ;Y7XW0aX/,a:ITL;/3>b4IW;E&Q^+KK3.G-Xc_gg<5.=T?.7b-;\]E9d
P1V4R)cLf6;ZQc29-EeZT-gY:U98V\WR;d8Tf3<T3#3<_N#17RGV_6BH\A[QV2A^
LSJL5((8Gfaa-=FdN&DI+;+BP?e46Z4.XPVDG[G,O;Z4\5fF[J\B3B2bgBf8@J&O
OO=B2aP^Y2.C;_TcLa=_:E,f-g/S&N]B;TA,\6\Mb=VRFVb;Agg^V5)]5?A-b)9&
X\E&)C#gceZ#-eBL)A([4XG#8)2N[7H_6(D(4>g43A0V[0T;WS=V,M-=U1g^f4Vb
8]C2&B.b?:]OZ1O4/)/4^R2L[BU=ZP,FH@U:MU:.,cVTZC92gW#E7KTYW-H=[(+_
4.Pg=NMTX#5\M@,W2+D7O3=JZ,.HcH0J>bQPUW+aN6FPUOQJ,&[2VR2[Y3+:CgQO
9Yb?Q.SQXg:[LL[TF_9_.Q)G_GA4(;3T(g?:D=231^=-S1[TZ.#E8NQbIL;:,JWc
VVgZU>bPQ9d@\C(//\;AUZNR2cUC\1NY?-KN7UJLdETSO.D[EX=.1aC9XL)_2IDP
=TGW.H=>C4E)@/V]Tb7ECJ<7MZLfJ#YLd3B9I#FEF&R7.+Q4eIFQ(Wf=8f.A@OJ0
cA^O02\bGH.\UD5G=M+H_](6Y.,;S5_K7@<Hc>;.3.82c-5U1[V;^F#+@SQb0^,)
<NgVb11KVc;S2]gX2C9-,J<2VBGB2-HbW?XfWO.,(/P]Ob@JZB6/\A5EQSQCV@/:
39XDNBBU/b)MdS>4,83bQ&=d1G1f><-J?gA+5dbG@:C6e&\aR:39aE-X,^#d>UAV
16ebc]AJ/UO_Z?,egPENCd>?U10&&1OAD7XC]aXD\aH6?.W6HYgD\G;OD12]G/1I
bMX,J@=?GT4\[7&KN^=+1-NCS(T.f<,T^;P<^SG:_>gE5PYDfa<[PebcFbY\GUT/
?\OU6:WTG6\F:TLA^4F5:\&98G2e[b(^W>.AEg/EU893798^@g8X0&W&-^Geag0L
AA78dR4B+:Z2FJUD/@&(QF,2MASeOKNE9GMVLP5J:IICNa>Q;O>_UK1d4cd-TCWS
[R&F->@]-][QcAUQDFb]#31R4?64NA+B+d+_7RFG4CPa2]e3Q\&N--176Tc^g_D4
7/+DS2ZCCMVD><&-(P^T=e>C8B2AGJ20a5/61e2Q.;gcHA[R;TbJ,A>SNP2(VPS^
5\(,0>3VN#0W(;f\S==C0<b\M+4F3d[Q@QJ[][e(6Y+#T0X(S5XbF#X8K.1<3WQW
3ce073f5fL-GMaQR/&;f(>M9:._H/3bC=UM//_L_8)OVeQ&-=A15eK^#57=LWaT7
NcVKL12N_\2fd?CZX1BcY_gVaE0(ENO1S^g&X_S0H-[6[Z&034@:7AE&5)Xb3Bg+
aWB;TcVgN)K#H,3H^Q7R2B_8P9#?NFB._7WPX&AG94>H,9+C#>PJ4Y>6_(ALcVSM
Ef[@?\A7#07)_.<@b@cVHdAUV7_?2E#8C#^K/#,f(XF/(O5Ra;bVQFV2;(cF#?9U
g.#8VZ?RBO=&42<@SKR59&W_:YGWbX/OS&;7YH[=T/WWD^@bXa,&JN]38^5,fZ>C
LC?+AU-\\P[#a-XMCE;W)QGEA-W?##(QZ_7caTCfTS\M:D:#REgPL;WB2#[V<]<c
51&7MeB=TTeW.7@7459=Le):@8))5B9QT8]-a9@BDNJ31\f)KDK,I=S<8,?B0BAA
+)_@S6/7W<F[(A4/KXP1/U^&T9ND\P9TPOJJ4QPe4TFQ-[9]SJ+fDNP(T6H2I=Sa
]K12+]?D]]gZ4<0^Z_T\3YQ.?dRA9^-[Y-_T4Vg:&CaA/6<aad<8Qb,fBMM1/D;=
<MfegE)eHc74<<V(0T_---?E&Z3F(C-F4BKU?=,ZK0Hd<)-aaB0[aS++Z1I,EP4M
g7.&=LOAf-M7fc)Y)>2P.Wa+DKM[>-:I7+Y4bIG5H44eH3A.R]6abR(+4S&/E#XL
(dEg/A/eP0UVNIe_-_^dF-/>1V@V(QL6-_B]=(]-UZO^TF_QM3ccB(+N4FW8]PRf
@cG#2]N7>0b&#TE6]^cE8#(7QdDc>:VUU(RX;U<WDS+9HFag5+_&gLgeAcM,N07[
_PN/6D\50VL^1E1aH0J[>_(8M)1Wd^5V?&):0U\:50=+dM#b=T#+4,TU#D.F^ZR;
MHX&4_2SG&:Saa2d-IQ>.>7bdU@Y>7eM[QBEVRNL.aW\K-B7a<O68&_POD@)0:VG
[)_7aebRW5=T4.6B4OA?ZXUPASRQB0+X9K]2OF#TKKX#JeNeV36)1[R?D3N>R&@L
gSW+_Ic;\1.1A,#K:&)6eQgS1E@[fYM:3?)G0c#KWOEW4PA]?bW4cdb^X(^f@@)B
C;a=L&d/[9Z0_ON[:7MX2#F.T80GP2DCQP&.CHb5@[g09/eKK-//3P9C?(8-^Q>#
.WAD_0e,6C.f/UY#;C^6(BX5DFV&C;@7_g56W^g.5V&cX+LA,7aC7(V32e[AA,M<
Z=\/I@A0&AL@>N?c5)gNU>UJdNe>X:+AJJR1#D<cUIO<BcZbe=5SU#Q^<HFUc+\4
=\,?f7[aO8(FR/T5<?a.?HU5NDBKf.=EUME=?5BYe2W-4>63WPA&/JdE?4^bVL,F
[4g2:(I,/4f&VO^J7=[IT\SUbTSg>:(:D.V1[NBWJ+U=3>J[c6fV8fH5@+@PP2Aa
,;2^>e7O01b\KZAGPEK)5?A.336^Xf]ff\M?[>>U\-C3a@G&;JV?DGKEda?QBP4b
3/#a</DcD<W-C^MVQ@_=M=#^H6=98bKbKdXN<aJ)Yfe8_=R@M/gZ9=RD)[BW7JUA
_O5L7XP:6]I>S?HL;,,;W[0:Ma>DJ,AgDA1?._0[1aV@cdCdH63OQ##2(W3Y,V&I
Y6]&IT-F#P/1d37,&O-M&R<>[SdSQUYg(&L&XVb)5.F^f[G+N+],1&f3.7b#X0X9
,NOYP^PO0D],]UcF2<LROI:+CdLcA(@+<4EaUUeOD;CgY<G(_b4-d+>Y,]Ld)[cL
/)eTBGR0IK3J2EMD9HUU/(7[52gR.UO_@W.J_SA4cZ[#VX_5GX-:U8O6YEAB(U[3
0_635Q<LZLWG8L)_/WHE5>c.B<-#+?bTN71I=_#;Z6N..F13a#U]f#N#bJaWc[S5
d<-X?Nf:02fW7&^&FA9OKaAa5fBG2QKU:C8IaG4A4)2[,Q)1YX]6H_M4[KQHGKBa
X&e:PU_G1X3(9gNX6?AXURMc\Y_AL8A5PST&P79>aI5aOUHdQT@;AL@@^63Vd5KX
5^&]>BZe3+V4:1[Q9+9E2E5U_C03?fU#e;b?90gT@JgeeILI]6\O3KQbQ)RWg,0&
bS.G0SV11a/.@ZgX]Aa3TLJ33f2)_,SV;/X2J7J]bH@;L;2\a=#BEgXV@V+/0O4d
X6Ca:QF8[25EYQJD>4LKf9U0?3O]5:2\/Qb@3MKa7PJLb9_eHKA.dbc5Qf)E/_1C
a)Q;.WY0Hfb#AdMfN^/)Ja9<JP[M)g5G7ZK5LG4\&DHT[(W&Va3UfQCe1-V=eW+B
>6L[0=N[09^KN^19BZ=:.XcTecK<:01R=&VVO=1Of+;IR+K_5K?9#W\HJ_[^K&4\
;IEB6<baDJ49@?GK((0F#S[N39G(fJTd=00-QU/KOC@B:.HK(JB1\@5+&\2d90cQ
1]SG(c,MQHGg2B60DT,gWR5#.BMGfS/>Dfb<_0,@.?#]f/K8X[\>PKO2YP]L75#7
G+5:190A4V@<R,LRWX#V^F+1LWOS./O_SE/)J+BF>54ZCPCLH@9C.>_W^H;\@(Gf
OFB05;ZbMb4/RS@#T4?MOV;GNQWUCCM@)U@d@:6V^bRSgC(3GfT;Gb/FD^ASQV;.
>H<WN;-1771?QfC&U)S2NZX(UZV#NgQ42F(+HAM).@S/0QFKb.HdG)-MNR5Cg)7R
GS^1U[&CMB#\SHN>\.84XgM)=:8Hd?YOT]D+VIB.D-68L:=,N6W06EK:;>BM1Z@I
P;[X<U3@#G@b:HWC(,EcIN_H]R#VH24f.Kc,_AFZGZ5Q<=RT5Y(3=B+b)QQVgc[C
1<TIa]:^M)=C>f;H=B?[bUNO#f-_69+Ud7eb;Q,B,-^I<-8#TV)U2E5/-9,082RH
CS+SI6\(F+=a)4V(T3N1@.0:I022JHc+4N.gc(3G8L>+0BTNYK6,G@RVPM,./_9T
GFd=:BUP(RgB(fL[a<12Fb]F[ROT/Q1W0,eA?][,#UTaBY+R)FW8bJL3_1Nf4&UW
Lg<\1Y)R?,JA5)fX5<CJA2();7IWTYL;O-_NQYZ^9-5C)eEe7(MQ9@BEgEFYER\6
?ISEKUGQ&_cbI:)C^=SNQU^=\Jg-XgYFcLI\>:R63CIW0MgQa8VZQ@5,74BSbL5(
64DO?;9gN+Tg)Mg9B6BS2LFBW8e9:a8fX5#4KRW[+<Y/\QBDd]d0fRLKG_AKgf0(
Q:SRGM3f2&BF)39Nc[bI5P6RF<<N.+EF:?7F02b7aCIM.W51)IK3G9S-M5.2WZ:7
FLOg\/?E-/5N>/9=HC6:EN0CR\?e/0,b)L1H(C@8;=9]-K5&5;b^3&^[XTXfD+bO
J(-:DR9CIe5fAbDGN-:F9U0EQ=@]OT1Ve]5/=1+&Y;9\H[_,#4;G3K9QLc\\;B6X
J5N;=a>;F95IBP[d)4D443OOU+Oe?GJ@;:J8Y&9S95KMBWP_BdX7cJY\>0BTW-V:
?.NSTG&4)Ac)R(S92g797_ZGGg8K0A6BCg)[_LKMeG0#BLCJ[FD,L[S)991II3TY
TI[.Jg5L/8/:^Zc&I6)\9-F9-8J/7D>W=dX]_)4HS_P602OO[V_?33c-+QSGSW?;
5M^F(\@TbI6UZIGf9KYQJKWEZA9@^?QYFCLgRAV^=fWKI<_bNARWS3&fa7KIHf5&
;1eVG(80D6HAYLC0YLF^KS7R/:9>-gS)[I2Ae1JUJIY&acJ2bCM.g;)&ggCY6fd.
MLDDQ\4;^C+3T^J1RM+A6bYI5[43ES.^+N,e>SbS.1b\1]@Td>ZYF>.95Uc0b8\(
4:SFL/\U+XS;>VfA,_HZ]DKGXBb8bDPN_<_C_QOJde-OI9e/DOS)eUUca.I8Qb+6
YRE0MN.bT+d5/=UHf8[F&G_CNA6@LL4K7Te<49-6]Z0f>\B)668WgS?fS7F@</X@
:V_4AeKFH@[DdLF[;XH30aTBXT_Q?O8PX21VFF1HSK+5/-8]Y5MU9T6K>&O]1WM4
PO_F;@)RcL.-Z8CNLI8+:8=aZ)aU(KDW_RQ-dMBDA1E,@[_fE:4O;3R[531\3dY^
CTT1U,FbT]EK>ffE/&)KZd8WY^GbVKSY\=D2Y_#NJWOC6)(8Ja=VFQW10.OU+P7-
.KVd[:FCaIbX?S\7FIX@aT=dW/U1J:?C7\V3RaTBGX32g,[WV#J.GD3bP0H+XA;Q
[(<(3-MYPT:_8GA6GgLDTNZbf3BL^TZ=<1:P2QL/B4-gB)\)R]D?6UJQe7F&#M?T
W9&QJ.ea@@VWQ>89S<)X\N?TVOEAVDANAU<X)e;UCIA,]C:GKAg_B8K.Df7&Q09\
DU^F0W&^=+MI[gVKF(7NHOD745+BFa=PS<I/.\M.W7a5?N71R[5<>[Z_?[YS,)D,
L1b-a8@caBVfa7GKCH&]-;H)4_S=55L7-]H(CWAM\;&FVe,2(8@a;4I]F@S/E,g^
4O9OM\<@bL-QBUDT+0HaWUT,JF>0&RCRJR1YGg#NWN]><9[LHDQGJE/V64JT<U_9
;d\&D1LKT>ZJ&TYf,]OLe4T2IVf_g[S1bO)B(ZDOQWW,,N7W75?59NX;JJ+D&)Y9
Y3ZL4YA[XC96?dZJ]I/Og2B?)N77YFM5dZgU7;g);T4JF:b06@^cY.9WJ8G==eW<
.W7=>Hc6)16@ZJVO/?K6bKb^2EVU85E?#6H)fZU//FGK+gH2+B1WB:6&^R&PGL=^
S1QP532:?bf[L#RC<H3T219BMQ\QI#Sa_UE:@cX-UCQZ0?f#?XK,_Z6=U@P03I=5
<K6\[)1fT]6Q=JON15MW8#36,4MK\D3:(J1A7<J3E.>P,83[A:[#+UJM)G)d#)D[
L.V2YY^fKT0FME.6TKY3;2YG7>/9)<GfP+\;_#DVD8\OadeYVK7TR;Y[0WIF_6R>
OcU>4.+MJP2.D#E.3a8?ccda^_U)+JAQES&OJ[]g;7I3<PN+N)XYf11,5..LL=8_
TLOS4#=F]4.E]N2S1I/0YP]S=PP>Z(aE.ZBaDX4C;e]gb+fT6YJ7P9d8Z\BGUQ3+
FO1]30Fc3=LPN<Re8SMIKa^^PJ33IR\UM.@7Z5S7dI1AbWF4H-++]D7/2?,LMXD.
]=??IFdX<&2WX>L37Y2efPaX^@&;D1<9Mg;T]2MAOO&)D\@bc_(#71Kd0A0<JGPf
gX2b8S]YA@W>MFP/8=3QT4fg>cJRF#H7VK=>S7H[>c/UNeZ(=F@[8a@U4<Ta=TaU
<ME;9WTdI;b=[[T@:3Ic[@N0L((ebFC>\FP<@R15@<>V>QD\=>TSG=)<=G^e>dQ)
2MbVT>J1.54DG_VGS3?XCWFMOP/0L_UOWeCPPeV)3Ec+P(7eGD8d[=0.ZYF]6]Z8
]S+&+a[5JO3?0FV@gN/.VBD)fcPGSF\ce(7Y([RGC;4D?C2\6&\[CK1)=C&(V3XP
2X-)A;cMQZJVe?><AH4?Y7aI1.^>O#aTRTg]B.7+(L&)fN)NJJ[=A6WBV1g&B+=G
Q5338)H=(/_1U]F-21XHZR.-I]V;+DeDQa\a)&5C<g,S&dE,.3=-5_f1V,_90Q_d
=B#@=/]E@K4+M#\1Lf:NU/[N\-/SUg+@UVZCK9b68M2DB;-ZM-VGC#FC@XA)F.Zc
.92(QLG/][b],6<D=ZD18gD#EI+WT/Cb[)6)c;R,NL>C1,54HZ4KXI[Cg2HQ:U2(
/5>VN)MM+Y.1P&73\,IFe3X,9K=c+E:]0:4cI^,SICP_J)X\2.^dRTIFca.[FQd2
fTR=4^5J>)V-Z[BgZIgC<;.GI,Lc26,SM;>H5b+7#IA\ADV>.FZ;51E4P+3]_P,+
ge/fCS(-c1R,4,F82S7gWOMGKO]O1KYgFFO8YZfB,Gd]aBOc2_51A4UB88:19M,W
NZSI)cC\+Za]KS<+e^PS4TRZ@&=).^SBWDd+52PW[d@D(]WF0-)fXbWaGCX=b\FW
@5V]XD3G:R5I=TUcMf[cQT.3A/T#;9Ga-CfFQ,\8PP7^<V?a^<R,D]ALSeYCLdaJ
]#BAG7dggQ21_YI1HFFBK2.3-5YTdAS4/^P2.WNH7)70;9(FRO<GFP-^c/K2#aI[
Z>Ae@ggX;91#bIOV]W]]-U9LZN3A=SW&=4d@d(:_bbY+e:@?9bf:Z;\42J;>INP<
5]Tb&GA40D^#N8.K^(@.Y8c?(>SE?dT_cGI1Q+@>H:88d;0#;L@e56cfB\cS.V,F
]G(A7?LPdY-NBP9<:E#bDE1#[2Y-C8<#_COE9/30=8#BR:94T<?SFLEJ-Q_6^V-8
gSI)HL+G\])>IGAdI:E(cD4[48VA4V;YFR#B2)/R7R&6I.0]HQPWWA4MDNE8.bMa
TfQ6G#KX;@e,H>-ZE3[\QJC@=dUKP(_V3<WMB>@R2USV(45:1V&S2,&0#e,d&WZL
/S[4ZX(_Uc(X;MaGbPB)3R)\?EI.gREBbaEE9_PZfXeXTOA3ZKJ37?0#341H>BKW
0a3Na@56;)[D1b:I1S_.^0RcOdK+_;Z:_;]^d2^aOT#R]DO/T4&O?9,>K74QKIgB
2AY2<\^/PHg6>.RJ)7,P9BD7NdL82K0DC<BW32PV/=5]9W:14/9CNaGXN+)cFX-_
CNPc7TK?EUX-<5-1:<ag&N/LT-L/M;16.9f1KIU7aK#-L,JCWfF5USC.ZD5YEcf>
Xb<UUMX5\d<6W)f&,V_=T7T7CCC+f[?LF9DB],O:;QP4?[bPJb?A^\Gd8ZQ]&aV_
QKd3M0H)SZV<aCW/[GgH#0,2;8LQZOEFc7]/Me=0/.OU\a=b<DFK=\HE[R#<Q;(c
W#e(Y<Hg023L&^QVKFTMVM[.X?P,B@MA[I6I07\W@56CY,)02c?aKf)9J+,&@&1K
g7SQRWC&LfUHM@+5DfggcX&)5\G,9U^Q^5M@^@)[gg>P]J2@MN=#6ddZ^D]OF+J+
a(^Q&D&.]>aHe.TC687(^OSN482GR=CS]L#=E.XI(_#TdYA&;Fg8aH/+G5:SUEaa
A9g9BGg2A-f-=)L6&Q)EV-83G)NMS1.S/\W439K8NS0K/=7\C)E<\=]B#6g2>[,8
QM1<QGL]F??eL-EgP&8Ga\)=A;B\U1c=M3:0U5fb-W?VV+D<0K0OB5;eRLY7;@5F
8?H4eGe@9/aA3P_RgbQ>)]8P[FE9.D7Z,:JWF[L6N=3@c^^?+W#-IQMH4K;,8^?W
<Z#]MAa2](TT=LJ?V8DLgFEUgKM[eLV5D##5Pa<O3C<?8B86)P?N7]6&J<AR>AQ<
(:b72MAg.V0MG=CLGM?/=\<USOR@G3:/?JIN7;bHO-[BFA31+,UX-DTS#-F]NG)Y
MfV8_ZF:^V_XB+6/SUD+.(g)(BN>;9?#NcL:4;VaHd[a:NM<)6>)\^PKSCTFNCB/
<Q<2[]302Y+,/J4=f__/7WUR\V7(:cJ-TN9?;[EEXC7Q2+9cceJM;6U#1&^&^E&@
D[)0X;Z<a_gT/bba/O7ZPbO]DWd[I&BHLfXP]K9&cLHL9Fd@CD<,9=64BD;U@FRW
7^;\aMU/ScS2]FWKABM>;,a+YgAEGdX0J3:<48cbUAX4-f;:^#fd#Xf<HFOU5O=B
&TDcI52O[aXP1aK=I)LJ]TTWKD?K+93eG]?D9#-97QafZL<:Q#66LD=PL9R0M/bA
5;6H&EX,F6@8FP(03SKVdHgBK?eOF89M=eJ>P>X\UX11RgL-b36Q+4-G:C4#_-KM
cQLSa20\[d?,Y1/ZPP4YKQ1)>6>N^eTWUS\+_[F9C5;^E;6:V#HL@F^dN9<<XGWV
&I_1\Ad:&5Adf#N75&17f9ADAQK2LfD)A-X/fF?R.Tg)-\ZBD(MFZ)@N5bGQ)2?Z
g,.Y<J^<cC[a74DdX))74B^1L^0bJ31TT<L6JB].MgT0X\c,5PHR8:b3c?J(<.PJ
+RGEKC>\;A)2<-^WL94,cZHbN]KG7&X.3Z(bOaC/6\dO@c&^e]F7[&CQOc/fVRTB
OGDGFH<L,-f:d<2738Y2=\J:I4?TB5EA7[aCT_#88S<dGE_1+;(J/JQE_-)8&bQ2
gD+a-;c,Y;b.)NfW4gQH+:K>D0644FO?8TR;3[(VM&\A8-Hag63MIbO,X(.,5K,_
-Q/K7VE.g:?80,>HH/X4E8-Q)3Z<8W#[@3K,,;,6R,gP@.-gUFJ?F[7WL660E8W\
K&P?H.FUQg=T/ZgK.[J[[:OJf;/OMX2E=Q0>#[FCLKD,KB:?6bD-+0_1B?7CX?2O
#T[=\X21:]<R5VR-M],bgAEH1T:8be><\GdTc<7G^[E06A2Q6,.F@O_DO.V.&.7M
K+._=0[FIFB)_4:FBdP8A<8I8f3&b?4Q<<4GfUHD#.2cEgLALG#ANJ7WbDGI=[(#
JCP.QV?3RSU/X7U6&;\b<[f..ZGeUBIT&&USEQ)K4UW4:IMFeF<>^P^BLb18P\[2
AR86c8,/_Mg\#4/22U5BO&RZ4BQ99G^M^D3#_MO45XQINHN^GT<7f^\,#Ig)JAUR
gXAP;eOOH-YQS3X1bH^fZC444;(cVJ9U1^WW7/ANd9+\RDX9Og7N,V&V9LdVA3:O
4a>WZ5W:/c[U-&OPNGHEbQg>MW[@_+,]>[9NA9Uf+>3f)]R#6T4/UK)gSJeG4IC0
O)QW-D6I@4;:Wb7@6?0aP7SdU,Z^3=PbdAT/:]/[.&P)8I#f#eKL\W;8S^_IYSJH
4cdY4_W&1EU9aG:@>B/-c=C/#(Z=_Q2.ae)eXgZX9;f2[Q(AX:f]ZCSDY5Q874D4
5H1W_@#J[-3D\&F3(PCPaKY-S@;\Q#PSS+6I#aHa?=)EJdf_)eXD]V^;/?Z+]Ma>
-^&;HZ[N&#]:F6AAZ1GdI,RB(cg.&P)J.M\f])@SA,+>F/8HXED@LH@<-0RHWa@<
KOC4MK0gNC9EDYCXH6b@JF>#/RPMOQ2E5a8Z>@.YN(2#=VXHO0+P;013BG=+CAH3
X;Bc&Ld3GQCD^0(FGQ-I^K\eQ2#\PX:J5eK6X9XL,_J69[UdEI4KQI1Y<2K5J[5J
48J3cBe(I2CRa[6X&^/9M8GKNc,BP=S1;W7RY5fB2Y)aa8f0JR?2K6NP@d^27K9U
g3]g+65<W-W-^H6W@D:ZQcCdCgUMDLF23_T23.L+UP-O@HW7)R5:OMd8g=D2<VAK
+)a32(A:HO<B.2HNc<B-P?PJ45\V/+G7,JD7eCfE8R\JMC0Nfg[GSA>X0N#V@F[O
>X;bfAI#F,K)#MZRV/c/+(T09M>^UCQ+Q7;H[B[-H@QBYSP7RVO>(,8SfbMF73UM
@DXa.=,g#);88bEPga5H>#,g\+aK]);_?_M^Qa\G[^EQD(3.B#P2^CXQ4^[YffWL
C+O0:0D1Bdf[\7IW6_414GB8AHM5eV&c=gS-c@9)gP==[.B)g)C\[;gP#(7>+\87
,DeY9^=##YG>[T61HNU7^K?(9C6D+K:_eR/=:DZ5?Ba5_@4Q.O)\ce#H,R-/f^Nc
1eJ7Q5CNQ2-eHRLR;JKf27cAf/c(;A]]ZP&7JGb^0@G=_(CDQ++HO>g@E^4:I91Y
/_MX5=9JD?DEeGZg[Qcg@8&V)45/LZ<V41;UT;^N@&MF:?PO\IdH.^gMMUN17I)e
0EOOc.;8+)D6U<7MfS5@G>=e8C;[\(YT27GQ>P(LJP:F8Q)UC14Wg3aUX_eBg1(c
J/?bfdV:R:N43;f:_Da@]4bfR&/L.fQVD4B-fg9E&D2F+4bG;PF#cQR,(Y.Y)5+<
\)f)K69E7Y/9VD0Je[a.)7X9?\HEb&_PN8WBVVU=a&Mg/Q3[\6.#1ZWJ4gVDO_.6
3=_[#<Se>#FB18f/bCY3..FZAE2RIBYS@(<J5gg#ZU>I7/DL2^^>2Nd;C0GY8&49
0:)d8Ef/H-D\eZ=VHNfD[7VWLPP5CGbJ@3MI+@e@aZF@IA6W#WVQ1RG8bcI<OH_5
P:WSRE>2g.WTV0?L4?:/NCR07LdP[I8c2@B70;]eGB/8_<I#BL2f#KO_Bg\LR4-<
J+c#?\3&8Z&&L4f,e5RG9J\0IMM)f/)79S)&#AJ#IS[XP=&U>fbAB69MEIKg[,L<
@cSQM2e2VV>^4@O&Wbf1KZ2&NFG4BgQ>@)SEFVG]NYPc^0(f6b1=3-EZ/J>L_d)?
_G3E&A<C]>&gd/0EcGGT=&9KM1B-?SaE/R4G+2;77fKLHP.OC?S@&^cc8VG\-6#D
)]fcfM0ZQ9aHf\1+^4Q7J@)09@#W5ID_,(H)4\?&4QgL5E#WY6&WZ.=J>FAMK@FR
ALI=+PZV#LcC8[@d6VAK&MB5c/BBdHB2Ng5A0YIA:5PO+=)D;1=GA57^JY^+7]G?
]H/fX3<>d(T\dY+_@U0E5-@.D-Bc705X)4JF:OX)@1K7981I:12XBQ&,;&g@c<^?
YL?M6-4aTS+B&eL=NMS6F:X9<L9DD)b;BJWQB?TROa+]AeBf9KHR:U9,&TV:g[_#
1W0MDN#OFb0^;9ddLeRJaY2&DEQ<H=&]9;/^,:Z5K5B2],#;OE,:]6K3)bL;9cTR
IT^JX>J)78UYd)ME&N9_-G0;T:SU+IHGD-4+=91f+Ef/ACQZB,4H7:D^:/_MDJa:
,SD3XNC8-;F=YTF<V:bJ5[0bCW.c.7IB[b3QC<+:Sba4SW_\-M;2)gLT]7g?Q)JO
O:3=W5Q9):DET(^2^#&0CHZYY)F/LRG_1/B]&P_0Q-Tg9e/(HS=RW\U_Y&@]E+Y5
FB0d33R/^bNUL3#J9C8E9-c8>G2V6NNA+I0@#<#R,YY/@S5d>].fe0>QC=_D<b(&
@2e_L7[ec?)a(,Q7A[1C_Z@-Q3[F^]3&?+W00eL;JbGNS&2Zb:@/#1H@=+G:3U90
b0Q,@cYIM=1OWPeT6?0H2PReYaL<PGKG]eJDHQK;X4WOK>>CG(Ze/+3VNWdHaCfJ
+G1dAW215M,6D@;C:>#JGaN]QVNE(TL:GHS-BFD7f.d0NeD;9]9HfHQF\-GFIF65
O1ZS3?1]H._/?[S:0+/9[JVc3R1HHe_c(KVQ&)JDYL.A:12E.OQBc&ML4OBUfU<D
e6[+7.c_gFc?M0RgX>/6)8I/Q>7F/36:ZaU;0470_/F9^-;64(@MXB=ESEH021RR
Y[P&4VX9BR8cSVDbWFD/EIXJ4;2+1Y1DN40X;DI5OeIXW.]c_4c:(6O[X>Y\7CZ&
R]>d3\(5R=?I48SH<dDBbHG@V/&afNY>],8#0-<cb1@&bT/g#Sg_XA,^9g@P4AK+
OS]#2L:.R?DIgB+<W-1CJ+)Gd(e@@NOc_S1#C1LDIc5_.eFQH5OK^3T6KR+BeQdJ
9(,]W6GJ5C,R+7O8b?g-;M_<K_OKd[#4>4<R,KaBC+)@3YC7[U-?;><>E2JWY83\
20e9D6C(E5Z5[,]fRDKOY2[2aPg^_/CP3_EOfJJ@<45JD+94UT^TORJS.,E)-)NR
R7,,H(?bFa=K;_aC&-S4f8B86^XRPQbEQ8S;aefT?IX:-d2N<<;NJ&/8J\e-[LfX
7#5ZN;-HVeYg(<&5Xf6.^-1)3^ZPE1dKPgcKbTU)dNKAF2#ZV1c=O]D@1S-dNM-R
27I2a>c5]F&aQA44;ND#ZH9(+aQT&e3?YSG[c3c1=CRMe-,3HS[G+80bN8f]C.X2
6Q-EH2=,C3=6PFS]VP>,=VNJ1d:#6[25K-6GK+_E0.\?<&fAO=ST<]=c5^9Yb][e
FOE-12+O4R>4Z&<72J5&[#YYeM\[Bf._I]a+gC.W095+eDJ,8+=.64d6Q52[-WPc
6@(5&^DW<U\DSA1,F]<K^?UCQW)0aJTX_b,B8/,[J>L2VgF1XP1ZbFPWELAIBZ@G
AB,>62&\&W@]U3IJ/DBL#Kb^S3>?7P<,C00?91NM(#dAO4a3-0=GcId560&6N18#
25>.37Lbf?X:FNeb4]^N9.)7+LDIV_50F9TODbS6bK3aFT/3d3215MeSHTR)WX]M
DELC=Ha@8NP4-S9^[I\LeATJW0?_L=>Vba<b-/c-b[Da/2JX/K+LP@4b9Y[C[D3:
6[R6I@N:Q<8-78.c8c[COTd4=@HEfWa2@QL-2>HF0@YBUcbTRYG=#CW5(YJDAKN@
\HW7b6e6()ce2^cF&:AVbA0d:H-HC=K<g@3JESB7B0=77K.F@BV.Af#AM8-/9BF,
854Zc.d>-C.R;]d[Og7/5_Z@Y6_]<2]ZX6Rb&(F^-N+[V?5<a(_d^6J47dMXccV6
05(7c5L)9]CDL/0<GO(=/f,7/=C,Bb4A1;[>L26U6dM5EXY]NN.6A4_#(@36:WI\
bHX_5WMQ4?+F1ED;V4>>-EbSB31P5#]f=B=@88+Y)@&P<=ffJ76B&G.6X7Rd=)-d
YMHO1Q]]fV\SaaN&XG)8bG2Td3,g/;cUWHR)QYR2b?KQU(c>MLBLR<HH,K06(M(a
)(C,8-KP-L8)J)QS/_fJ<0(8Q,bX[3WX4ZP97PDW9UbJT4caQ<SO(AGJXbQ-=(Wd
;P[NGIaYHR]8JK3_>5V^O^Ae51-Q=9W6P4-0\H/^PRSOE[#\H&+OCXQ/A+^W;G)[
NL0;PT#Sd<L&L:,OFJ7d1e.(@CW^Zg=1Fc)2SW@@2bCIE3X-5N<H,^QTG<f@S:)9
[#;);I;&?-;;)A@Y<Pd)P6D^QBK1CQ9GO(9E1f?NDEACUNFK)GHcEcSGD><#a=@K
OI.\[/?<92JAH35<WQfXRMI3>[F9Q/0+YcA].)A[-U>R@]e^B0[1EB;c5eQcNS/=
305g?8)D@\14C^fV6aNQ:)8g]#]K2TELB5e\c_&UPSVS12Lf_Z&<B.:FY::X4^48
0_&A4@g<@1^4=J,c-H.T8US@0Q^J@C#YeNeNNC,Y=g:JA68)aF&UMReZIgN6LLVI
L[7FUBAKJQLSA_d@7RRag)Y78=10E,K^LeAAQ60Y1eUBeV,G7BEH0,_2)&OJJ,^T
&CL0J/IY_Y7PM0BMWLQ:C8RaMSZ?R+\F2?XJ+a2MM;(:\28Nf[SH[?9Z66E>f:#>
-QPSCL_5ODI+:[/Tg>E-/I;]<L17L&5@Q38cLZJ8FD#)6#)\;K[3^Kf=.bN=/?W>
8><<(B>13]L7/Z6fL?SdAIDJ1b1NUeg77SeAg_??##CT5eG;4EgWMVLIL_OQEMP#
FD3Lee4UI-<(ZOP+Z38,@Cc/&59+[fHMX)KR=\O2EWB5d85-(4I.Y0E6d5#8OEIS
#F<=G41@E(B^=5,1V^^90_2.R13G/:^<D/)1feT:;)>V;5[+4B707NT9F>dXFP1W
HMTMdIYB)b\QVTZVSV3RB;PXPN9Wa[BgO??dX,5<?6QZU[0Y8KbI=G4A(1;A:>1^
-AS/6;bdK#9W323?>XeBRc[Lbg:030>QG)W4/H4>VI4IQ;GV:0Lg7(@ZI81@G\G8
gPO_Z()-gLcFY_1447[_5#GZ)ICW(OGLD(1T<+D8J.7IRS9I>b50\PT<LcWOC_V+
5HV(G01c.\=&_/,FY66+9,Uc5dAR_[6U<&<c)0RabH)_0<)#I90d;HD8?&+L.#2L
CJaNX0#dU<N+7V]1gD1#K\TV+P4;74__RTG&7;10_8XKCePZ+Y<N(.ggYQWT6XgU
1/(dT[ab;5S=OfV0GeLF:g+TD_/FN>c4HTXJcQ?KgSP<=fXUWb[ZgG1@R-8CR2(g
X)f8=f1d_79^Rc0&-]3eB>AdQ</?OOa,(2bV976294(6G(DHgIPB#QV__,2Q_9cE
aH6?)HebJV?,=?77,3EAQE^_(b,BB,-\E63OfJd>XFP<==YCWSRc>@8^=0d,;RR0
CHD.WW>4Q+\IM.(\\BI9cD8+Y9CM\,M+;B8D#L9Y@_Te1+QOI20CO7V/<)NFS#:K
T\be,HN/#06B@K)/BWdJELaVAZ44):fe/O._F?EOA,,SPH14V30\+@=C/:^6OW;]
;9aTK308PQ83;PM>[R-D7a7=dE3(aGA.<;HaNTY0W<L<ZRB[dZ<IO4116,?c&48a
VSQ+>S=Fb3H+Pd]G#\)dR=/cAH/^,B-YM@<0TaMU(=e\6=5M?0VD4;YYAU_PU/I3
^;PV-G6#IEMO?.c?EL<W77=<MGH](CF-a0bXO+/6<INB0J&I&K;MD?@<G+P+,P0f
R@HIDgKYgcVL[^G#NZ@)[9J#.DD-Bd6SPa;-ZI3g(H[W^TGe>GDH1OISdc)]M[I;
Rc>aW0RdD.J-(4/W4H-Q(D\X+65MZXA0(V;[A<5XZUb,?2A<7e:_f/4NWUS9E?b^
E@&=_EBO6+.#6U?297CB2B(Z-Z.0MX>Cg712^1T.DE/\]^K?[N3Na0)9LJDMWKaD
L.?YDVG(,f?7Q951#/>-3L]20>;0_H8aO_6Y1Z80e\BNW[E_;<H+HBEG4BWL:d7^
b]^Wd]JP^_18FJ5fISbARLEdY2gRB+-N;I;RP[J-DML;FVa9#<>)D+]@LgBCZMS-
H_J<K-9R6QMU&ff@X&fRdee\92<,d)0U3dKU(Z4130?0^^<JBX;>WZGdM2>#1SXD
]I8FM,YX)[8\]570Sf>J&1U?N<8;C&3&COgPSYDP:74QQFgcLG89B+g2Gfgb@[^_
K3DEP@;[&]Y+g+TBBAI4QL&eG#E&4>S8BZY^@D7Ya#5355<Z_V@+C^9Vg,M5dD@2
-5:<b_^]W_4@NIK<@5PdgB:,?eFP5aDFI>?^6N(F46eHe-MN84E7E^GE^1a]ZaRZ
;LQX>\[OK.9=NG([:MY\Y(,N7bZS(/_9NT@;IR)#(bTdC:IXUR1SPDUg9TTb/>I/
#=U0WL5+\VdO<V5ZSAK)#Q4&;#DPPM,@fWGC4S2KL72_V8)H?4@[:(C6>aD75G7L
I_BWQVW807BW9-BMM_LS96bW?,gV1eL)+4LIE6R@bBNH?_0U@VUeO@,/__6gAFI.
#g31>\XQC;X/-1_RFCJ2R1c3?<N&RGELBL,0\5T1?.O6D=RQBYIeQ/]F6UNf&B4D
UbR0=DNe:L\ZP(+6RS8a:;N,Z4Q976eeZKc36<=eSXIQM9BK.f:HGJ#J6d=K-6PG
6,1\+DY0;LKgJE2dSV<f^)&F<JZV]1ALg2L]RgM6?g.K<_.&SY:0?f48&Z2L@ZII
eLc@.&I\bgEcfX&cdH]F[4(KK39V1\APEY102Q]g07FP@bHNVecYJbD)=3^K^SQL
W>GZS5?T)U1&EN_&E:VC;K;7.IB]S9;Abg:JXK#Z-UC#Ybg[._#Ce,cRB&O@7e]B
]\]0(>VGP:EO3R:AM839MU,BOT0XY]HP<#ac>PFH@CHX8]O[=(,\P9bXLGgB_ABQ
Y?F#)(^g.?7Cg:SN)Z90<:@+728J<4#DI.;B<c+b_CH80<<dHL[OW/(cC6(-g0bR
e#HMNF@W,b9//30\3.-4@))Bf;>-VX>A]O8VUK\+KWY00#BC(fX0+XW.(MPgSV1g
TDW7CA)EP:?>BF+L=C_MH?9P5egf@4<eG.f2?Z6S.R1,K=\E^SB4&d8)gY:XPZ6<
@PcA2X4@L98KQFegU+,&6<gf9R28..0Z)aLKf[^bf3SM\.#EZZ,Pefc:&La57Y/T
>gSUX@8N/FXgK]K:+Ea.e8e&;+G@MBO0Le/3U#:^bX)X.L(_9RDMQ#E8S,6]aQUa
,HO2OS-cBK.OK?T>7/=QXNX#g]Ng<89OUHB4D3a8a)<F@8N6,,EV_^eLYSR8MM+R
F)X-WBPG#b;?EaD[.^B-I48e04\(.QD?IL\SPM:K:BHYRgGVMMPUN^0GDI=G^RbJ
V:668ad7(?24C^+T-EG+?TCFFCOBN8e[2ZGc+8Y/TQG_FC4Sf,&G.I(2L<1FFQWO
4ON/O8\D^R/EeN4V@F2#-H5151g#?3O=1<TY>WPFSBPc:P-0J,MOc8cYR#8578YT
C;/0d+E_[+/RVFBZPD(>?G0(3)6C_F(3G+)&2[[F;U_G^aZ45:F1+W8<D;d?5A_2
Lb1?)3AKCc6O[4W?+V#<.@&#f16:B=6W?#a/We,<<d-@&a8BNf04]J8JL#21BVZ0
0+>[CH[]b8>24g-]/).RD)4GA],Yb7HQOFB+F<WG7IVUJ:>(T>[)KPWf?[(U=?.A
e&/6QDGV\_/20PA^PTP/=M9U7Ng.=O1AC^d+&@B7?aNb.-f8dGMB<b5C^_T04>91
>0cV.80>?LO<Gd6c/]22g0/A;:Z7feB2N=MAgZ(,;SIf6Q<&1cC+2g]UBW9(FC-e
+6Cgd^PB75dU8G:IBQJD<U7C+]8XE\X>/X+@J<&:NfSJISIN<&d0BO4E^Y5L2dP\
>)QYeAaL(?9P@a)8/9+QS):QLKb#H(HPRDe?X(gMc)&.-IGg,AFgOcQbY5,fH:M8
b)C>/-2A:3D2YQ0H49G6MeLdKH@dMI.a==bEJ+(_(V^7e[^Tbg@-EBYUT\_<Be7W
>eR6QaZa(c@6#FffMUR5FI=S.-[YDIIaL[)KaLG?0:B>/.4[9#?E1YOBFY6O(=Z=
dC[LOM_D]8?g\0&fG#J24:LeIcU+SP:BXeMdOcO=V93GBF>f]6,NcJN1/a52EYF?
c4#bA+B(\4Kf8Y]Y\19::64;T#/\<8#4;AL54#>HWaUZ]Hcd+O<G6T<@[c6Cb28?
Eg>/G3GSN?B0&:W=3fPJ2?\NFVV\Q-NXSX8U\NFE_;d(=0CVBe)AK.Rb0P^.#+:M
CK;_D<\XN1@XVV1aY8_O9UD;FS^S6=.TA\V]/,:,+;a_?MRMP9EP^B]C6F1K=3BI
c\B)T]A3^c+#J=835,;;5ddK+aCCde>X#__:^bcH^ESU5[X8VO1L3[e-3A^Z(6SA
6GK=QS/,82C.F/NbXT?[EA@_cJbd-:&7W[_,f.)Ja?)NEKeX]SE:LGS)@.:1K[fe
#RRV+AYJ\U8XK1PTX1)#JZZ;S:9NcFLIDVY@YT0T\F#>W2@]Nb#)D?A(Kb@bYDG9
<N1:)Q8199HYcg-ETL\.DU9\>^?LRdc8_>]bFe?UK_N?AI5HeAAFZ80P4NLAY=b=
TP\\D+gTbSaCH3TDf_>UX9M&SALN/X)O,WJ)a7c1:?NIe7c-TW.TQ@1SJ6MSdC8<
@UFDg3#R51580U^^[E5GdZ+A\+(82DJbB8R,;?Sbc9Y_d@Dac8e;2#2]?0C:bdc,
aN9c[-J9FcO9V5GP^(b66G&3b744,gY@_(1.1HJ>)@-YVET87<E40(36XC=._^NN
=0R-V+KG&92Y4geNaEEbe,RNNe:(aO1XCPWfJR&bRQD1PM/Q+(M.fdSG0O(L(Q,6
V[D#8^7PQM]5&dc0#9W[.\-<fU=?LI/[.FBPNH3\WDV(^+FHE?>U#F7XNRDI9\dL
TgLa^\0K#?,[F:RJK;6a#<dZQ#OILBV#TGMWW-UFTc]#/2IG&dFAGF^8]HXQd402
5U\2gH>cCXG;U_@B9X]2;-P])L^VZPI(+WRPPIEPDE</;SC72;],WBV00ZZa#IMC
O3),V>)a7Y)_ZCZVGFCTJ0<EcZ(B16;)0^Z\\V;[(K(d[V0g_X:a92C6X3-M:XN7
PH&E=8^(Z8:-@#0P,6/);GPLg&:^-/KQQQ>O^K6]DfTQ&+Wf9<G_>]S3[S2c]e1;
f34T0D1T-VPEcMHKO;PMK+CEX#cK4TF_>2QW\=Z1.7NE,TaWN#:bFBS21/2TIL)G
C9G:YJXHf,]J[JgUQF0(3JI(53dNNVK@J_?Z):#10-:9:M:XdFC)Z9GG@(&J:OMC
R1[ANX)WHc;a\\RD[SI0-&4PO#c?9=5-7<Vg/AK92^#2[_T400]C5Z^Z;R7Rf?#[
f8(7[Z]GgVSAOM.KD4#)\:[)Dgg8XYPBJF0a)Z^Ib<J9O:4#D,AQ88+HaC]72eJb
U2UJf34)I/QFTa>\KeX&d;33,df7Z4fW3[G@fL+9Ed0(??0H_TNeGCLO^Gb3VcNL
CZ67@AH0/B&Vd<Q=V>1)7+9Nba:=B5=OY\d/^.^.=f6J&J3a3a<T>=,3N,O]PLJ?
A\\)55JAWX/T-_Ba4::(PG<V<^Xcd1BRKZITE7E2/4UUGDcbWGWD#d;bb3_79=g>
\d,;^DJ?-,c.c,48M+&L9fZW0@]WOZP1]eGKT8c=U?#/3ObMJ>)U4)61/>dR#DFO
6N@U_V_:X>IE<4D.\((c#-D\O9^WQfD>#,b97QY:6+1BIZ],+W@e45Z:-fBTTK/2
J,IF/\<ND4.8?FgY]1e1^.2+D@L7#,V&@U[(:3/VI(T(J80TDG1?V);I?Ie>6O7<
=<0:QK&IA[,G,_7._V:G\GP-W6^-fHgQQcZcSd5WK0IW[d<gf>>M14MNHcI]0V>G
Ad9H5BV+PW^O[LgB[/&AE)B#bfb&8Ja\4F4[.G(=M5G_^#GbP[;M^df.4ZM^OOAC
Y+#E3c\9)&GUB27DgMbO?6d0=28Ub_cK^)8\9;NRfF0Z+IbB]][4XNM,aWXE&2.c
4MYHdO\CR(@A--QC7Ad[(@]:X_a16A(#C;</Y7EC,+gS;()O7VFTIK7HedBYcHTD
7EI6EEZJD_@@X->:9c)QN+.C@N[IB(FG:QV6Q#=@Ta@.c[5L&?e&_&@_F.J#V?DF
,T1=1=&5T96=2/Ig:Gb+4OM+/=SFQ?U/&/2H)C9KEZK(I6>^C2H?DE@d9g9/Bb#?
N742=_fY;1NWa/4+_[H@_IF74a-UPQJ2b3?@I&dQ^IT5(IIP?M/,O=^6RJ2V05bc
GK3(EXKI]=Wc^J;LH4-a)PGJSNFd/@VQ.SJ/f:6]7dEVF4J&RT_BWU?^4AK4-27e
Q#N#>5=PG/68P):48LX0.1G(DUG^c0^Z^Q>L#Q8+N+QMLFAU]]V]U9?3g#H.3@EI
#.^,U)7U=+&I:,^)8.dA+,P4EJ6_PI^WUcO+@J\8Z0dSFM\4,)c6YV5e#-g4_8cc
..9a(\<;1SMY9I<G)48Y4g:[#M^FMg5X#4Z3.^P@Je4TMUEHOYGOf^F5(,92L\,Q
SKa+-5CTJQ>#7[9BcKRL\,S[,H3-=NT_4LQQGV8H0gGSC=IeK;IfZB[(IO&:.24Z
PJDFY0a4\>6&e4b_c^R#,4c^SI_VNDgSRJGLfM7bZOcWO6C0[^AcWB.\a_9HY\#)
ZBCfb:M>)[&QR/16Ua.?gR9<#)YFVL.AddcALOcN+N&=aA[DEZY8RNIHR(Oeg^C>
0&];4X+[0@\:2J<S-Q95f=9e+@S9eS?[+O.cWR.BH[3Qc_EM<WLFOC\<FP[J/5[V
RS(L(\AA5X0:ZeC):I3Z5@@F=G+#MPH17E1BZ>dN9)eGSE4@0cXe,V14EdW-2Z](
(-4W;RKV:.=L8OH]Q[6BE28S;6S#JX+R19I0Y&/GEdM=9)]=(WMUC3XRSZdRNQ(B
K935EB0<b37;OR:P?3/-f#TOC+B;fcJdA[AX8Q6_C<F8QV>JJKNT/b<8VXcSRLXY
P\?a8Z40=?=G_IT2ZA;KED5:_HZV<@.V/+\\N+-]=d32RI-8TQESO[P+\RMMg2Ve
fedNdZNR[)RG1HZL-J?<]IIR4&V,UKKBZ8P=4KgdFD^059gggEM1H_3/Ia\f,YS#
R3N[A_^CDf-Be@X&L439=e+EZ4VL>ff-_U^D_CV0Je(JV6AP<IIVFH8^4:;\=9V-
1(&6_K+D[=N739P:OB&B2/_37,GOLLG8TWe_Y&K[AD>)?:\PL^dVe/]/?b.[CA7\
e5Ua+F+@aXP2P]CM)IM3#3W3;[KN:L58A,-5UGDa43eJ@;QS589f)bWd\0[.[.S8
NI2.)YUX)H[GQ:Zc]+44M3&Q4Hf_BG0D-,K,Q8-?/Z1<N<4&aK6N=MI_C1N0GEJ+
M>E@&-[J__5T,Od^bQ/GJ5I<0UM7M8[_f0JP5=8fQ&YWX:52fN8g.;ZY-5JJ,H2R
H^,2.PgMM=U2?((V-&Ma<3.dVbQ#CPY:\(I&ZfgOfNP;L-,QeGTDY,^Eg8G_?<-5
ZS3#@68)8\]M_U1UC]XACJXPEH[=F.VQS9VP25O+?4Z+9gM><g4J;JL.UE;^&OUU
b07]f;]4eVNQ6?HJ7e(;HDU+[?TSAIE>O7,YVA]U,MJPO)NXV?dPJVSF?HZA5&;V
b[4LU3G5gJ<MS@c<L^L/7,:0b@SQ4:C,g\DR<FYUD^H\#(U\TO?9PD&<E^:7.P:G
+\[3\9U:6B>^1aa3TG_4ZM)[2S^Q7baJ,P:>;,Z7-)4:JQQ.MB32FX10-X@CGH>A
RAD(V><aIK[PA#dQX7/LH<ADKaf(eb@&e96+WH_1PU,2e=(I,L:Tg<]S6fT3L7KY
Q^b5WBR<5V5=80J\YF\NL7UV4Z-7:gHPeA9_(ZB]bLZGZbc8/04.5\NMY6?=2SaJ
0@DZK.,dO0eXNd#;TSAM>f(cHRY(6a/g&Q^U#[INXOfCEAcDc,bLb;)e?#=H5gc3
V77>A4)VUI_LTK_+69<->#]Ze0OB&.OXK+E/6>G;&;[B<INU_88fOcG_REgc94\H
MYA46RVbX7-Rc[1D:^QPaW.O#d<N.N=RdfGZJ-Sg:8R?(?^_T/[RXNTcI_3(4:3e
G>VIF.d,L\<57NFd)YEU]ZXUR^Oe=,)VD0ZdDDeF\7aRF>OSB8#<R.U.^^HDf>R\
Z@HXRH5M>HR[1Re>&COPH?Z]@3MH^Y/AV/^O2GgR@YFA.NV(=@4)58a6@Oe(BZL#
<=#-cR3QCaG6g@,B;/,P__&5JM-98B4LU,#GPLXV>[+eK2^6\:T8H=U:M7U]3>><
b5#S&Xg@e==8^4:E4_V@Se[=_EQV@:+C&W4#bgYPVgV82]EdBIbOK0D_.(9=HdP[
LKB_-c+2]]8Y1\&J:faIHUTc>3PP7cTe]F.>CS1\V=ceXU=[]#eIBc/e4c@7)OH=
?bXCTc]5.7c\MUJBO]Q+#.FQ^aT7_B,F0+_,#?7X>ZJNLZ(b?IO5E4\-eMCB]c_D
DQKKP4)MOJA;=R-+T7F(R[DS134XWe(?D.R.&YdfG\:^N/c3@UPWeOSTOZf\N/KZ
0)5LI96d+Q@Y)#8>IXeIR]J)-YIE0E.c2_XE4)G=K;cO9..QR=^[QN;g@>>PC=_]
_-39K<0(;DA>>g^Y=d@gL/b=<B(387DAKb6Q+Z^1HK4f0386f_-5_g499#J-M1IV
WBL[3:A//\M6ND[:c8c[g-KODMS8B_)V.K)d?116JNB36#0A5\YXd<@LQO74PN1F
)S5U[EG,QF\?dNX349+?fKCYQ&U^6fWNJ2a9P(?(.KA)f(TJJSRYJABcAB7U.TK?
QN6KK7QYQ^(J73)fZ&gKO+4FOU;_Cf+eJGdJd,9,Q3^X<C)>P4I(O]Cd3IL=MOB3
L<1Ib(R)JdG5//3bBJ5@9K@Ce/BVXdI?I3a(S1G?OS_CBa,U1I/egeJLIfV:J#RI
<<#ae4\]bZT1Mde?E\NTWa=F5,)8(/SF/CUGB<&6QE>0g?SgVRH0f>J4ES>CTGfT
C3PbDN\&)^JBG>gZa_\b<&3X:MTJg8)LJST,O+S=AA#1BL2Fc>d9EIXMA@:;]I:,
LV&AZD\QNW4NY6@R/bBJ[1,\X6Q\0C8.AT\LJ-KPY^WULNSSNRa+&B6#(,&AE&RB
:(^MVcQ[D,CCMccN:CQ4(=,X?P4<Q.9Wae+J>8+0c88V:AOW^OF-S=W#7QGOd_EL
>6&+6MRB>=QW+8ZUOe+#/5Q^9_=2/3N2S:I>9Ud0:C>_fFVATV>+?-3:2MGAHR\I
[B+S(6LOZMK5aWM>6aa,A#KG:::];f3-W?,M.:>O/XQfccb2CA]:<dTP]-16@GBK
\T?F;^QN@73Y/g\3E=-Z;gV]/0#Z)3/7TR,25b97E^KaDJY6f.(_8aTD_-Y3#/A_
TPRYPON;BIFAbSIb)/6c#0L[67Cd#AGRTcYbJ[+_/GR5O3&MVP==77H^T?VA\a8P
/XbN7V2W0B2-D1)b57dX_PX<T]La(ZH;VXDMKKUV;/5Jg\c4=6P^ZJ<Meb.a7/[O
PN4<^2AA12+2GA&_-AWf1AYRd@FU[8-,I:/?^O:?/)HR+]>M4&+51I-dX<E]2Y[R
XZb)U=5Q;>61@#W@I,bM&BeY.c7\B79GG5[E5f/?^N(TCQ5_U1086EB:U-^(8U0B
=DC3U-=63K>UAOeO>#e9NW25#T(;QK@O@6,.PRGaDT#Y7gS^:K+->OP)/_BW^@_E
5XI45/C;M6,LKO[BK7[R][0ZY&I.;L+Z&?d5#>68@S^CBe_1\aQ4=Ug6;W4-.5Kf
]?PYTQNE_^D-.;@:7A4QJ:W5c&,RUf_cF1,PZ;DDd2d.:1?>;4f-3+OgQ;=33T(I
LH\X:E7X=F5]2@5PWF8>b?Vc?;Je#W9b&1\8Da?[KDP]NOP2>GY4:]ePf_gDN:cK
]@9?[MOI1NT4:KRRQIULQ3+fFU:6EN2IF@9Ugd+HIc&0ZWHGUbGdOe?]O?.SA#bI
#=0\MB9Cb<2.W?f=FF;/MEFTM0/WdRe29I4M>SB56.IC:P)6K#0MP4)-Q6_P.CY6
HJf..8J\P7#f9/L\]:G-1P8]-TWS2/g>cQ2MFFZ:7YcT[Y8-S^W)+XT;>FE888XY
_T:(3=][d04A5KKVKR1]#ZO3cgWaa#dg_+><W.W<#\81H@U<.R=Ib\B&]=0#-fN<
.O>ccM/gQ?E[f)LP]T=1JINIB>SZ./W,M4TG@+7-JOH-T##FJZVd:_M>=Q;P,[Y<
T-eH>_\>)?@,LR&4.OA80K-d3_@g=DE95<D>VF6dXX.RM6NBXP1;OIJ+_.bANT1]
M_.8@>X&b]HKc9O5G\S\P^CC+Vfa_a/_WE3ASI061T_5DI)Te4&CD_/3DEZMI--f
[K.cJ:#.TWX7KME<O\CfMHVL\?DRK^15JUDN5H5F<Bb))6Q3;J&_X3HU)_TeaHCI
Q>/;[R)QAVG,dRd)1.:B[R;Y>[(Y?bbX68.JCRZRHDg^V@_/&fc4W5.V>_&#)CRF
\,Z5Z8&L#Z_d.<-5,67X&ZRXOV4G#LF7HDbPXX,:B>KOPX;[N@K]:e[fC[DLLT_^
T+Y2KA,4T3RP#+K^>M>O.9E#b2J:=A4Q^N9D>.BFL1O;+PW9^;.^RME3:>bH2Icc
>1I>&CHgHgBbB9S\?\ed,Y<36)CO,+ZZ8_M1KVX@Yb[c]L.?d:+K\==Cg+c@+&)/
g=9@QcXYXdXB)^>E]]O.b@,,94YaQ]1):8b]6Y=[Y1/CIK91MeJ2MRa\0]JZ<EBB
_SUG0^(c^#85,X-Y,M9P>gAGL+;Ve<MT6#-1IWU80^Be=[.YeM&<63C->P/LEebH
P0Z.EV1RT/c=B&g:S>;-?/-/,(&(B6;,J24#N6E?eM[f29eDAV;g##A/3W[O6#Pg
B>>DL794WcR^IZ&(E&?Kf7>Mf^4R92H.-6<?+0aA]cU6JaWdW\2Cb4AG&BAN;g:Q
]C<0+O)QcMf4\(24,Ue3L_Kf0+9Xc^V.(AbC?&_,@0V6X514Dg;eXKcUJ1JE+AX^
/.3^G+fAO5K(=KV>7:-ReM6\+:&g[HO\Ug8#QJC+#27P_3+a^a[a+9RH?1Y-XfWD
)HU.3S&JZQ8BDT>]1>P_I]?/R9?L9KW<VU,E^(IUKKH81H1g9^.6=KF.7;1+(/]V
K6U\A4+E.C952AE0-7YSS1K6[I9K:JfCUOH\:#?LV4Tc-XKG_<P)MB>>#)QKc&],
WC#JK+]-P-::8[_fg&E53Z,JFD@8fcSMK.\IAc#Q_aB_:VIB@b4LY3@7<4&RJH.L
QHYK?/=STg](SEKc41Q<+P;<2:cE->8H9bZU(DE^9B+NCB@4AOD\M9(b(H,?N;Zb
;N)LBcI>ORENIb_c3=CYI3V3>beWa#YK_R3e)_P;YJWJA^C#03<fd:>OcJ0.Rf:\
Q:XY:0+AKG9>XU&B,(-3-F#-fQ3E>6JZG)]5(3+B2KQUadMF#BC2@9]g\c=2@/@U
X[&I6V-4QR,<+J15EcaU_L1dI]X[]5PO;D/faG=8_ZJBB3FN]OSLG7?VYJ_+XKIX
[CLAJU-RPM.de+27g4,.&0T\\gJO1c+:X0RP6feW42SP\S,_bE6:(A[B#4d;RdND
P(Z&IFc\A_OcO7LL5E91=+OBVMR;;dF0fV5F(#ZFM:B7d=LRCJ7TFK#>RG2DQ/?4
b)RLR9aJbeJg.;LAPNMfdIT.aVOE,?4e)^J^)a_LKb4K=T3MH<.\TIQP(9-]38)L
6dEAA#d=FLA0\GfM(581;_GJDXc7RWaOX8DUg6[a+N+6>1C;d43C#e;g)HS)W-(:
W\2[.J-<eF^NY4e#+K(I98Q6CgcPMSC1G#TNJ[#A+1IPU=AL^6PJGUD>L8-._ZHJ
e:VGKMMR340gH7K->RQcCVYFARaKB1EQ4;E;WBg1,MAJgTO<D>4#F#Ha/^GT^]:X
<YZ@EbL?Z43TeTTK;3Y^+=-KaH)V8&,4)fBSU06LgJL6W2c7e]1dKbSCH1SJ;1#7
R;YKgfI,F-O[/<6Sc@G@EAG;CCcbXB0]W/<6G5\b,.V&HH]QNgGXOOa^S\OABK20
eGLD[).-4,T.c1cVN_70aab&DYcU./#Z[9[N,S7&;:LM\AYPa7^ARb?g]+5SKZ^V
P]SP]L0>a.-TFGI@>U?6@TRYeKZ]2P31Y:b?IM\F8,<AIJDcP,?a+8+bTT85c^1:
4LDY-E10V;3>YY82,e[MMWMUaP+WQW#J]&?Fg(/+MFV^4JIVA8b^9.R4T(GGG5X&
PLRc.f.K3Q+\GPHR56IN^LB?F;ecC28HTRUT3fKXVTVT03Je];1&eE:0DNF75gJX
OG/8-IXd^dV5]c.E=;NES:&;\1S-5+U[a-eL+R4Z70TeA-)<M>1@gUUO7L1H^IML
->Q;?F,Sb>aa1cLa1?(/VPd./f5U^/P4e6QTSORaD(eDXV05Pa[OaKJ_XK#EGCad
(?&I)YQ<Ke=Jd+-2?KcL)]J+9O##gT9N,LW:>a4II[@C\0a&KfFL?P[1:]c9<+U=
eT>JPJBZB]TQ+,EEb]cZgT;AV83M8>5H;RE[.U[?OgaC\^5V7(-HI2RBPL_T?(G3
:c=_6a0H]UdE(DCY;cGP72c<QXDFYM]PRcb^L&R\ZT8<D1I@45?038ZL9c&EX@=_
W^R^W<M=e@H^fO#f,/aXH03(TV[>aK84[QEYgI&OJ1C[6[ZRE>U6>>/JVIJZ-]?T
_/5+(-3Y\03F>>TS:P71931PMD((&dT[QWE07/VLcHfI-2/c^M:/FEf2:f:]_<[@
TY5QPc,WG3dARE49aFf[BLPd3MIYKY)HAA03Z<3R640U@G1M]^,(^a.[>&,>KW42
YS0A7?/\(Z91L+<TNS_V3U:+F?.W&=aANA^0H.UV?J3]0C<BW5&gLFZ3+]+LeaK=
L+1;<S]9FC3:;/a?8\A]F6cfG-Zc4ROS9\3TT=Y[/P#KHaIBFXbY=UH[MKZ>&;7?
W)#&.^D6CQ?Tb\Ld?cDDJ9PHd9J5>g7d6+F.V:KXNF]ANA<NP.OYD<fbO223A+]d
CZPUGF&&2f#Q@,f#X6JL3R23NcI[VZOURP:0a(51HF6.PaPG+.Q<Z-KW4&PRe9\S
BY(I5J95/A//HbD(2^YD??C,[C>BM0BZRJS#A\6#N)RD1)d&J]eAgXda;NV8_S#+
#JbVb_Ia[;d<MSQ,-/&V?)8K1fJ3>S-gBP^:4XR]\D5/J11U_W<8YaB8[[1>IYFg
SC9eUOU3S;IbQN3S)-S_B:CR@PO:#V=7&A[RN,PY;98,<aGfP:5OESLJ<6\ILH,6
E2g/(.CIRSeKBPU^3/+Vf)2gFZYHLb3a+<8638?2:?]_S-]+R):4SD2)5_/#>>2X
:bJ(VX-6^1[_TH5>SN/N,N#Q(B.P65Y9KLFEG>]L-Q;G:6PSG.G:4()W>Sc63dE#
N6>cXD<V^XgD]_S;BN\TJ,,]38X#e#H/RTdYE)@45-e@3K?&0#CRL57B,&\VH-U4
\[G7VG03)2INFC@EbP=dX6L]faU)eCMF@b<SNeF@C9AV8E7^cGL?I7W\(+;7J7gg
>Ld&5QY<<5Mf+@+1&&>UVNG?;X&DaELf-#EcAS7RdZK;@cZC7e,?FYf+g^49a(b3
f^Gc)ED(2(>:=?I@0+@3>4^7(8F59IO:H-#Q4;6A8eNb=:=:gBF.5A^\,^fT\)>b
X^=6XHg&C3#M&GT_JCfHIFdd#7SH6,VS/D\eCJQf[3AA2IZ4;,KZ(-=@/ABK\??^
\A6OST#G_9N8MeC\3)^C43[C<=(f2?H&>?@#8bdYFM^5M6[OYN\M.9U1,(P0_S-1
N@^F7M?U7_]5f[D_ER0ID<H&>7SV283,ET6.cAf,S+4cg.VIQa_COSe/S]:ea)+g
bUSH);g\<:_#\YX\2H7ePgBK,LPFZ1Q>5IFDE]1#DdM#HXUY_:N)G76&CABLJ@O7
B/&@MQYfKeH76?HYXONe=?IAfZ1H.,S:OZ<[#XR9@)D<bFWg:-RDYdYg\U1^_W(U
(b6b&6.@ZCe..P#HJ1,6[E1PA\+ZUSG(aV18PAN&6[d?d9(4_]:e/fR@G>KL6bAP
6Y@Jd[)0+(<(337gZ3+QD6Q<eF>-U.<U4=U@=8^?NQA,5[D;P-XJSGgE..@Md._D
^,E8>P@(ZO#&VO(XEE(7\0(e<US#;GFVGYfFW#J?,<CQCWE4a8Af1P1H1#NSB/_O
RXT4S2X?eM(ZXFdIKRMW2CW;3M>_PAbT;=K[UBK1Q&1?:1&Y8KSVd[LB8^HHR4-=
ZM,.D(;TIB6dPc1VO(@e9FMZebB0Kb+CG/FFQ3V0Z5:2AKfd:GcV&AV.#[fg&RD/
7fQX4Ec=X]5H@Y4GVREAUO_Jb:+J<Md4.&:;B<\.BGWHdB[?GPRJJBT86Sg8be=5
76b[dA7\905ZT6]-K0ZFJOU5ZE5]:g@]\08ZX:Yb@Q,e&DWI>90CDBdT0[6d<6YM
_)R.;Q5(+(G:6N0]8J0@R\dLJ-PO<<VWP+D=Y)HQc;Wc,YHeDc97eZP#W=KaS1C2
+HXRK064)T6?)f(FS:>f>@2.B\-<6[[PERJ7cM)fWU\Y52GNC#J\Kg#OV^9HEf4Z
A=D6)f;e7=85_O2-VIAD>9_/G7_3OPN\-1^H2O.L>EQf:B9YNMM:4SJ9U^c_>LQR
]U.1I+TDO&L[F-P?ERBC(a;X(@DgCKF<OWBTDBPSKda(_L5#f=A]aH66\3)YO-F/
6)O12Y7JLGI;]L2>c@ZDN<7<Y[fDZIF>?cZZ(]7bf5)<;Z(;FOZVI_QR1-16g7;Q
/(Z<S+X^eb,_8SJLAN[Y2gZ,]8\eKLI39C(]Dg,T&YH-(HUg<Z@SN3##7#1Ce;aD
H)OA0NK6:;)F@fL:cF8@I86_YC-]c?.YR@U8)>WGCS>/0bKWUZf-.U#J?IEB@gZA
ME2,9f#b.)UF9^X@KCGN.])Hf;7Q-Sc19N4YK;53;.AR#<CKR/LNE\e>Pe0\a0FI
]NHWR;c1^1[2;D_.0M&,J5df7B:Kd6^I3J9?_:==;HF6]R^e\#F^3gYgdga]#3>g
3;fN7(_U<94^bEX:a1/VW&E.UNZ1_?A_4@8FVLK3])POG21HgfYabKRS<G4I&?F/
-=5.NO^Y8/PMWPSKTEa23//6]74eNPHY^I9M:EgY&9<EJ<_cAC:A[MQT:\K\TcOA
C3L4G\f/e/L4>L9;XH=CQV.MG7&-1\WH-+6NR,>3)=&+b<=V3SV@4Ef;A]26:BAZ
.6a_\-OW>6c\XE>WRI\1Q=YJS8^)/ZYSd56Fa5D/O&UH3(UMCCE;)+LUDEOggg^&
6a13Ld21[/6E^F-RLR?\c+<=LR>gK5)G_6A?L0WUY-4JR1PG[72#2F)U&;SdB637
<O)LgXa,G(ffZN(2+gD5^G:LR115HM6b./0VOS=b6UF0(@^Fc^HOG.bd]V2>]FWB
3?HX6a/O_K.c.6RUaRAJ^K2I+eK.=-LI+Kg8_Y:S_B=CLc_[ML&=ZPP5K\O8(G3?
Y@g_,[+[]<]gdS<&\LF;edeb6X8WIE:OZ>/5R6\Zba;]]>;aKTY_L6G\bGa13/\9
]94[EA,,YgdZ<314e>V@4:9K@d(GTCaCKFf(8;U?g#(dERGR_UV+3@LKXPM<41=V
2=-N#<(bGGCc/B8?cI]?^K<YJ_5b[H=V]-gT#V-f<\<_a.QU1=_8e.b7>#).4Y6e
4NS_F:M[#YS7CNRTBV>5C:7ZGb<\e;XF)ED)NBC1<N8P6c&U1U16(U\A7>e2J5-S
ISITKg<W^GSCPW2^RV^]E6]^JFV,(22WZZLgK>_@55CbGBJ;PZfKI[0b?PU(+YJL
,DcJOR>LEJCHfVW=20>=],;,]T.G)+:\)HR9/=?IQHE1+6_LfXE3.EGZ^08+]+JF
V84-]8M8V7e[/=YBP1)GQB8(gM=6d2ed:Qc0.2:0)Eb^ZQCS[>e;NND4MUK[G1;[
\97_8L/g9[4dF-fDb\:29<-E=P.Q<P3V/=f;@gDWI:+NbY]E&a17eMH,cP24<3#-
CI:@GX2/5VV;JG5[Sfg)S=B?6gK=Z_ESI<8@a)(>AOggLb0N@G_.PBe\L3M3U52B
->KT7]c+M+7->H.aU)08&0>U)T,M8^M>B?:Q3QLdf=OL=c&<Paf0<4K73[Z=^4)e
13]7e..M=-_VUBM[\D[+-/N;fPOUQXc8=I[S#C@cQW196JLDd&>^b;N=M?2QZR+[
SM?0>cO=OSP@Qc<+beaOF0/&+B<E<0B)L^dZgD-WL6NS.?T\U+=_g(b/1[STC+_\
AF3Qb#1H[+2;\Le<:EP[?Xcfg+/ea/2#U8C7-B.MN8:U;:BbdAI@Q/B1=6>Q-?BI
VW8RZX-ceMHIP7[[Wb[eZH16O2;_/SM/a7O+DBf\LgaM1G;7]&]M4=[JO-JHA=MN
)^Qg^.;/0P(+VT^b8R59R8@WYf_.X(J#7b8YDVB#QG=_U19;:PA-)DCKM:Ke8W(\
JgP0<g[,JITd1S=5((UIP+c-UI^/4ZHOH4fUS?GB[H6WI1?O2I4:CP<3[KV_(04b
EaBg1dY@dYdaG88=XFP-&=Hc0]c@)FMFXR6CR+bd=N;9FY._T+/)9-HP[&BYG?,9
+\CNTDb4<CN@K;.@2M.2BXB(Mc4Ic2e,=[=BBG-WFY_/(/<S+b2/(BbG0e2@;U9M
-AW@.bU<D&;B;6Q,E/BAV9TaL=M\V8&GO-VeB#Dc<N05FY?5-2=?+YO@X6DP?+[=
5SMB32ec_KK=7eb?T^VKUT^TH)M9^O,9<[0]G7SI#.X@ZC)#ZE.ET[S<,bDCEPba
X?_0P]QT):UKL\(<7LYQ2[A)@UE>LXI12g?He0[1;Y#RELUceX0:7ad@S2/4_3M<
+.d?\GT=A5,dKY.[]^+KON\aY+<Bd&BE:\)3=Q4C+OYfCI076Z&:C0-1=;E0+QVU
9[:TU\0EDJOTUJ?^D__,9TFLPM_S7Nf#L5?Z2bf]f0].K4S:7^>X9@QB\]LWc[G8
K^X@Q&R,G/.(:bR>E,T(=bI99?fa-/eN[8U]b.LB\b-7Q588L?;VD<eROf2U4>;8
.P6gU3D2;2M@\eg,?J;FD@4LQC?#;I)XCW/VFK7I0VFNeZQI8J<>9BPbV^G\WPV7
cZRJ>^JYfb7IcA0NW+#@/0]KB0R,P6-;+G_&@_.Wa4BaEJ.aJ-=9\:c8,Cd_O\G,
>O(cWPTd)+#TcgQ#?9M0W-ZG6<>GR6K@P=AN+f/C,Kb\LIeX:)/A2FYGNd0?9M(?
F\YZVTEB0cL-AcY6C^,3_\X<Yg-KU+RXK_X?CW]g[[>W)IGV9W&A<?XGcS-.#8gQ
<&I5BbNN:Rd3\L78GGF0P&)33-TZ=#G)Y\)TZ\:&CYc);0EFEP@#4NM93.ZZbBNg
,g.2:L1?E8+,GBXUPTAcT0/7OW=-S2ZH__g8F:-cEV_J>9Yb0K&E]5F<:_,F:4:L
2(FfYBdUB^7M,C)H;eD1+^RW#1L..P/c^BBH#>&.X40f,DO^8XM)G4=\Lge4;F]Y
C,c,<d0WK,\e35:V227g.]9>B?1=\&SXO)]fAZa^=S-\bgPR]I3cPX-fMgJRPeO4
JMMg?7F-5(+94g7=8+M/_>,SEb1B8>_98CIYa\&H=,E(>Q64^)^U0&1#EPB@HeAQ
f<<X)@QLG<CZJfK\&Zg/W,;=H:H[Bb]<_EVLM+Z:9cFDb<AU&ga18Ac4]W7gF:0d
@6Q<?a]:0J[=YRDc/bQRP?cE+.EUV;&^:Hf<-E/P;&OIBW]AX8CAPHG^DBTAa+OH
9DNfWZMGfSIVK@,6/3VQ^Ie3^<CLN,DTZ(0cN\fbT<<P7bTcCc:b[\aDCC<_[VN+
</cfdAdL[d8=6aHMUPR2E60)IIeTNgJ\Z5&3(VOOO6T1.+a2YEd2@):89c:1a)/C
Kcd]0a/3WC[GMZ,f&#:2K77M(DZ_5RJ9Fb3?ODC+S/R]UP[]VVA&+K8]1Mc^<_XT
KUGPDHf_N1</6&542-<d_[^f^AAgXN&JKG>)9/^_f=IW-RJP7T&eXZ=Ec7^>c-:]
#73;I:^J]L5T&Ag9G]d^8O5(a7>TgfCSU5-ePFgI6&dZ)[GF@ab7d8_(bG^?26>@
2eED9.ef-:.L3UW)ZM/IS:eJ_NE#LfT29KHaH3B#,J?L0>0Ec5YTQ>bFSXd^]W_K
V=#TTOSI4-dCG@E?+c5A8L)>[=cg_G/TDGd>AAW++8;L1T[S)18.=4G:^<KLGRW8
aWQ?GJ1ODNAN1S\BRZ#Ocd[F7ILR44aVM?R5FJCYf+9EgKdK[B[WN^CK8d;4&XST
?cO/[G]&:\GWQD,^^;HY2(ffL2C_)A0bd+K_E-MVPH@6f,LXf)+IK:dN4Oba.QBe
4XUWecGfC@=O3Sd^#6da6^Mg@P#^#L9\(N]<X,2gJZ9e5Z0f(P#2Ac<Y#YRH^@9+
/63@AFb=6LX:[6LbCaC]AcK+d)TSA4QI;:d<T3GMdUcKQ+-fZeX?3#V30=)STG.V
UE0a))MF((&.a0G#@&CPKd#:gU2.[UA<_ZG_V_X4NM1S]VdDg&U?,M(cSFeGMg,=
L].???aF4.;LCG56cTB=fK6;LJbfEg/e#-bCVY0OE@_KHe)aDHd\Re3@cb/-BJ.-
ff&F)-a/NY(P</+@;\P3C=IcZU9@K-=4:;L266[R;HEaXOf&,OZ?]G.]VA-V?UT6
K3>7+=:;M,N;5dQ@>W/<bfIWQeCK_QPG?gH/+H#TM,3GNZcgRB+F01K(T,2(0f.?
4[TaXF;5Jc+WW@[7dOX&fL:A5@f&7a\.WVde_>PEa)/061P<>HecN@HCCS9CO\dJ
9NI3&Hf.fM=3R;P4:6.-OGJbA[?_N#KKC8#.WGI].9_;1fIROgWdCXI)2JYP4TJW
JRLN2>dC32Ea.0S[9M=RCdA#]J8-DF;Y[N-PN@Y5HcXJ#BPNF#0,dSQY8^3;I>,H
X8;H6d-Ma/L3V(Fb\d/)#-4VYRb?D\VEW7gO0f>CO0-G_OY(ag_>,\?1IKD[O/>=
0DcIL@[D2Z^T<,HfF7:W&QVB0_aGd<dg]U87GIO;R+NBY;5G9bK5=P;fZ-NdSFE5
/-Zb-:<\83Hc[@ZAQX6<B/gG4g?U,63@Pgd6^@UDILXD[E?gHL(#0=DRXC9<d6a_
4Q&DZ#NYB1GHLA2FTV\3RD=KWA9[HWZXPNfR;[GRKFVU,/P;;P:-\E_QV&3/b,Da
S#][)7a5A<<QbBHcRI4I__MT8JBUS<V>]<bSfa8:03b_1Og+T#0&/[J12\Dc7:fZ
c9[S4J<QWF?I6]JVO81]&LeSFXg16>7+]UMKDW^g^I9B[)X^O;EIK(YI<-03G[_(
I<J/c0&MROc+XX=K6GbV+80e.F#,\WQ2+WaI^gX2=&>,XH9bY;6&7,,eD9A0(GcV
6(RAW.5VN/YZeJ]XTTcWB&T9@#LW^N;V?eE95CQ5;PO#^[7YILO+I#Ef)1O>3#g_
_KQ4>@&d)3b34U?+Tgf&\TZ5399[V@[23SgXY5HW7S]KB-W1BRSLe>WU?KBZ@Ffe
2eUCMI;N(/HMgS,PHCF4Ye0>bFe=MQHE&^X,Y1ZJMJPab(DSb/KA&H?.,4<U_5Y(
H[f:eQNd&3bHMS;.:LZ)3/a8L;MV9_Z/VU.L)a>I^2PT(&&L8,[XAX5[=7M7_faI
(7e@1BWQb[<?I>g#9K#4##BUSJKLbB]0Z/>T61f#cU,=T,SOLcC00AGe8U1[,KM[
PC[,1-U:0cBS8UGPL508UccI2_CXB.I)6+GL0Ae)d62OPXL:dOXEI=<bJaL^VXM&
dB2X\KY=WP,C=Q8+Z)?ZWJA@g\b7R:&gcIA?(D=_9PI>=VK1BBaRR;bU-&\\A]dS
eZN[NE,\gU:<b?\YfTUL/-c8C.,@.MZ+4.gLf?,XQ2ba6eGK#B(5WE:[@@7N0[6)
WLS,1.+?VfW@3;WM=aa?MTf>aF>9P,;BC>;H0P061cEB0#>/WU9AX@5O/A0VDJ3T
W2-Z^?)H@5[A):=6eP9M9(EaVZeL^?fCD2]B2=NIC3d@;X(aR#>>,5+7cd.CF7W[
+2D3[AAK:YD8XJfZW_#I(0Ya3NB>KGZCPEL-8?EO:BZ;Y_<7]N_PX0E=^c_Y;OY[
;Z-PQZ,L[Z7<M8YgY)_MJb#GB&cJ^\R,^>aDaAMQQ86CdOX-<NVBf6>W--VFb-_4
-gQU()#COPQ;>@]F</B^XP]IX=X4-W1YE)_^&)]dc<b4[2cAcG3I[K(V_[dJF^8S
,A=C)M8Cd-4)PH/[0[a]:BCUR4FELGO)M&#B2G=P+Q.;3A,.5FT4RVELJ1SS9&8#
=B,IM[2S_b1.:a50g6?ULW)9H6_cEWf67UgK^E&RULMX7#MfSSV;4GRX[DN@39Kb
SRbJF6[,?G-SK5._aGA26234)V-/YCN9,ZdJQJFg;G=(HdKOKG170_K+MEKWC6F,
H-/Z&G&D:DVee[)6Led#DNb5Z0MR;=KW&Aa4)Hc?JfH7ZJ.ZF\^Wg>\:/_>eO>Y<
c@4K_VCY#OIIP@W)##<:V_6A;=5:S9fK+K?^@>X4R^K9A^[=HcB22IE&Me+C5+2<
e>G/?O:TbIGd3RG8(KD04R.]?>3Z<ZMS#=14fHO?^F.3X8cHA5P.O.-0cd8b2DW#
]ccTd[fcbU@MA+[)6MW@b8]84CDH@)3]fE_6>3BRL&7OCR9IIacAf0VHV1M7CHSS
a,BM6b.fF+CEeX>5&Rf]R.5(()c?2JD+XLJC[U/R0<\AJZ7T2,OD3V]>32;WWWM3
U<)GUa+[f>L?<DC>TXfMCFdK0VQe@AN1F5GQZ+HKIdB4J/3:MgI(V0Sd[WY?CB2.
<84.F.^6=KJW.\]>7M)ZXYfR@]>8a>6=61P[0UB5aVYIVO9UT[@cR\abL[O0+8aH
-(:)#(G^@Ka7U(?1(FcPd4<B/48X8:\;S:1??PP@SDJ-P7-\291;8f2=FUI&;3Rf
ea)@E5Y2HVA.aD:F;2TU59J.4I[9UKc-+SLJ__RMc+cc5f#[PKE1Z_\?>Z,3O5^g
ES@0#^Y]7@\eX1K2DC^NFMLY<ELTe<JPXcG#<+MSST5DZg.Jc-&0)C)GE(Y[^6,K
@5T?7Sg.>D<5RMe>>aO3B9IgPc1gb=(HW5AI<+LP;AZ\R6NfSB#=^)1WaZ/g?T94
5,\\0&<a6JXa2Q[c44-;9GCM<O<QV?RJZ4bQ(-9KA,M5U+:B7R(V#N5UcfUW:D^f
S6BQ9#S\g(>?DIZ3f@g/QbC:Z9FfBC1\LKW[?gS&-0NF)7FRIF#b#HA3HNE7bdc/
?5JJbf)G3K+:<:&=9Ya+#T)WKQZSC)O,KK7#0;_a;#IH+@[P3=3,:M[NY.BW8AF5
QF<08c(MOVUJe0;CfL-ROK&H?cO.^,>((C4(VVIDYH9(N_P6[,99#=_U/YAeCR-K
g+>)#8cJ>Y#H8fcb#,IID7Q591)_5gdKK=eKLbN4])W2/GYUZAI.XeCWfCgWPB>)
:,,N,adG^37\CQ(O&8:N][:6a78.@^HESA6,&AXT0P740MLB:HE^<,4<J7A>=8LO
&]\.ACXJAC)<]_(Te+I/E6-JVWXO+<<N578T984E@_OXH=DgHc39^Ye-2.X2\REQ
34JXcf>L?)SN?(\W^.2aE5-C4=^PGYOEK4@Y<8HFM@R,K:g;8J>GCCA;AX/QAdD>
aIVU;GJZ(b[/?M<T/X7RUSY8SN9]E:G&P5Vba6b6KG(f-KDN(Cb?#91T5b?=SX42
G;fF)5-+A.\Z4O(Cf.K7>c.\]49ZS4OCbX477=[2QA5D>f3e?OVRZ?MIPZNNWEG[
B3OD26[2=AVQ7Q3DUF,S]Z66B&+M8^NTWZ&_Wbb5+dB+T-24f4?-,K8B\AV]>J;.
).Xd]47[I>UE(66GaM-ZQf==KLc:?,]H&J-;@RHe_TRMKdF4J&H.Hb><3FTgA[V1
MSa)4Q#\-W810f:UWO]0\8(VgAaeKR1+>A;aRGB2CX/\fG]N,bM8TR5#/#Ee@Y#E
Q9fY+IQO1_,;LDX9M#8.Q.,8\?\1a:>+\][8^O_a)aB;E&SWCY^cCLN+V=S;#53W
a[1M_Z[c/d[9f=WB3C.NdZ?e,:f7N:(6Y9D/dUgM^b.eP?GfD(H0dGTf.Ra9[V#4
JRSaHf2<M+-ASN^<WAPP3;^3,U9P)80A\F<[R&+\LfX0^B@?^(?DRbTZ<V)bB4&T
WLJ(1?]K)W7gNggK:O+KbNcgE<1<V./Y1VB_R&7P]E_7.,A[U/9>(,;.f>Dd8/#3
aLBaLDc&M^Ma#a8NK50Z+G/g-6f=BO@+_[G?fZ<QXgZL(P(=F3Wb:NbR[)Id_aTF
Q.d<@[\X[>2T8Afd3HRYQY6L[,?Z47dI7Rc@.NEfVYBZ6c=ce=7TB_]P&N6d[9g7
K>20CH4W?IZZNU01GW)OePX\\f50Mg\A8K+NN_HD_.N<7\G,<6YP1+)-g1[OQ60H
)\E\+ZMScJ<9F\H2=H.[SH)dW::Z:A?g(OLXVbc#KKcK1A)>Nc8)_F8e1afQJgBQ
+GU7Hb)RIHD3^PU<63XUN=dAf026?RWg3cP<6^V4U<IdQ;UN5#?TM+@FBJW@I4@M
-SeVLW(e/8BLSH.d]4^96.?=U9=b+X4>f^IA?#g/G2YXK+.ZXUW_+\7X^FL;@#/B
.D?c_S2e8dYI7g9Vd8).X7]F67bNB)OF:P;BJN?J1F2_:@I&Ld2FG.LL@NO9,9Ue
D@<W-._LZH6R^T3WM/Q)4c+L[bKGFEA3=NM1=2)DU/RQTAXVV+L5P0?F.7,G0?.5
@-F<-TK_DMP1OLXWUU&gGXEQUIYG<SHZLYN=EVFBAN0IORdTQWc_56M?M=9.&VHP
F2c)GVFD\RHZ<S\0J(aR\WA2@cd9OD03N^JJ5-[N6@g0,a1g\<NK;3-<SJW\RR7<
03Ze1d^PS?e7ST&>W#BZC.A\(MYe0)[(^V30eb^dVgKZ\I;d+V[QY>eUWP87<,54
MK&RReCGOaU.1[cNCQ&HE<XX/6.R5]Q/<2;RBf+4f>9[5IS6_d5&VS^,JcLa.f1?
>H[D:d:(aY;9FeGA,7<Z2+fJQB_cS]gXATa\K_P_R#7M<bY45O3G#A#TN9X>M7MV
^-?9N7>2Z>P:)-#A(b]NKUGANS__,1ZR66fKcQTFcG#MX^GSDW+N^fQO)T()B06b
SJZRWOZ0b4XSB)^HeaXR6HF\bF#:VL&,bdS:@_?0L?:=4fV9N)#E9_b^AEC1^.XO
KN:TU;[c/g6b2.LK/3e()A4H-[JT7fMP<&+TCb)6cA7#79#g_W<8.G)D;>e/G@4?
Q5=J\-EQeV[60C^&>W>1d&=D@d^K//7?(7:(deY0R2PYUH/VMW#B4+S&7:Qc0a,Z
QOI1S^F\QU.7+Z9[;AP:E2e+YFIeWRZE5S-XEd&(JF-[?3CJFK^4L_.8[1HX0cJ7
:OVC2LW&\EW;VdC_WN6Q0F+)b#@]Xb0-QS>(I3]ES9Y4B6\PR8DY3HBL)/QCd56e
da].O#bJcA<U@EUa<<\7d:YRbSPE<V[WL[[fKW7M];]aCMGLSS3O1d2SCV7M>4OM
Q#XEVEBF(>dK^V)=8,MMc9)5+TTP63CMDFIX-dYMb_.0A/f,f2BC5fJeUd5fEG;Q
USRaSb]GWNeCQ>+ZeIDaZK4e5[CUG6]?Qb_Ca>d))Ig(fO:)4?>IA;/V2X/S6;d9
EY#_7IcXJ2=91Z;F><WJ@L=PBdR[NQXN#^gF#M(g3J-/ZcR=7dXM?#N.>+[F-<9]
a7,J[)fY\c=)YVS&-#=4DT4#W,N4HLCC5(?5e968MIa?7:dTW,NENdH<_8ES1XL2
OCdPG]IH]c48P_fD^(B,,e[WIVVeADA#QGR6/YfK\:<gT2&:XY-@fFe,=gQD@:1?
7OeadcY-E)3.SY31_@c4.&c;T;_V5a5cXd4M1,(3CcSVZHOHYQO5E5NJF8Y5ETK.
HdJS](g8:I<aWe.<TLM<&fFDI.XD0XFW)D^f].d&?LGX@cJ?#3TYSG-JY:H,.10Q
g;/=?YgcXR4e8@:I;K1/()Aa6E1KfCSTM)YS4c](>F>203;1C5YUD0RIS=W9<2TJ
C[Q=F<DEW@L>VC9&)AO[[-+0Y\42Y7dP;ED2a&^@aW8)EA>?+&D8<FE1e=<:a0DL
)a>eYR&.3cRP^,JB?f=\3T[@^9NS\>JZRB[a2:[V_;42X<DLXM;SDMI#+QMPY4,L
#f8aLH^U[5JfSb0bBbXdH:Kf3D;A8=1.Z>FPQ>SY>T0GHY3e72?a5,GS+d-9<P1&
+]OG#?:aId;,FL(Q3:OOJ&OJ/:@Ad9P-PVD>L;f5<F/?OFNPd.aD4fU?0R-65dCL
>_7+Qb(^1gf6W8PCg0aXLAN57^3O-].U:(e+JZ46PEX>7N(2RP;LA+V9B2X+fPNf
d6aGAOCM3PT69g5#8,]d&H:HKATTK:NGX@<[Sc6ZbcVd^TTKc[T(XXV0A/-T?6]K
dfL0[:R-0)P0FI#;M#)HcMU_J0:)[7@W_d;ae\AZ#eWR,&JA5;XNPGIXfM&]\UI^
bD1\.IS1V41D1+SE28gb1W;:c[;J[9?^XT(\07PUCJ/@+SNd16@f+LFJ00I:#F#V
-<bI?a<#DQ7^g+-aWYB^GUL]Mg?eK5>.K@8PP10@OAO[^K))K^XQ[-W&gH&L&HSS
QV55UE:Me-C=.A.645gQL-@QF2X.\gR[L3\7ZJWTXV;bZ#/R7gNeR_/[aNeLW3(<
A#Q^Ue;T(#B2RS:&1ST&RE3^bJMVNS/N+E<ac)2M=?UWT>/)a\6Y3aCC#TV?BaTL
)GBEJDL.,]8cE9,LKQ?MdYDV0_E?Kf@LdO&7@6J,OeGFXLP&./H,MQ0QaY]]OX-d
g:-A3WdM:;P)_.:=0eW,D5@&?SdQWVA@R:W@(F7FE[8?gV=]Z&)e=8EL/6A<5YT/
ICC\G4cNO[,.e^/)W5cNc@HJR>-6MVF/I7P#);??Y_a\30R[K82dUQ8g3_-F]O#e
)T.8/4QRH^X=^V;4?07eXDA._RbSEB+2ZS?W)f].K0]MOX^NRO<.?IQJ(>J8U:LS
e)MU+/KDR5Lc38-HVA[<_;XFL<I;=V9#XcBIQ0:d8L@7:b\Y/3Jb9f?]K_bR68:2
_GV>;)108&PRCb,BQ\UN^#I1DDC,;P1P&\5;9BQZYC5APQC-g@ZXP7UV]3ZDbb_/
6K(3_RUSL+TET&]6]?PXPaQ4dQf(XGHMRFPGKb[(2Le&<>-/b[f1:B+DaFG+C/\;
;b;BBBLQ/EW#DZYc<)8UX94.0g?e>Q=eA([g&,Q+S_.^XeQ4LRR.&I4c2;^MgJ\;
R@\]D:);aD9D.g.X69:gcMP7/,DCNP9YLLH(O441Y6H2EbOQID)&<_OEA5Tg11F0
(@Q#7N3F18e6P&MZ4>OG7fTgL\7&?+PK>9Ha#@938NX<f]XO?^<Lf#&3,e1dD/=F
7gbK.##M,+W;2=.N)&;FV3gQXN0TAR?87a=.cUc9B-f=&KMTW-cT2,9a,&VLT,MI
476@(EPOX:/D/MgS-@[gX?N)?a=PFIN[Hd18;\E&B<06RXJX\HGT.IQ]Q#Cf\,Q;
/#Y52_,DG(0-YU]6Z&_-fL2)dT@Uf2KA.P/CLgOP9EW_Y\]LQ5>&R#NMIL:K(f[M
=+I#S5,#EfQbYg0;,G7U,\<LA,K#/JgeF44):fFMZ\F,GC.&:;]6P-Lgf5OMPN-0
[g9R5_+\@MZ5S6dP,LPK\.B^6S#0#.?gF1Qf-fUG169=B)/Fe:5VZVd20X(.Y(gP
O<MW-3J_H@I.5]b-R<4?\d#I(O?gC+2MacTRD,UC@e;-T_X+fKYf#SJYB[c:f^f1
7WGX91W-7=5[1:8F=SYD.4[13.Ib(:W_M<N/gNIUCS#0RR5d1,R].aFL_+b73P-f
]#<DXTI0LU,\(F&P:FP2Y:#X.88\>dgfD=9OM=3,RD:C+GSKAJbJ.fZAX_2?-[H]
Z-EU5M=:TL>eTXA)WP,0\J9HQBWNfI57.Z;4#GY=1H<FRH7d@(5G0f\e8PO&?G4=
LR7V^afSA]:CdWHCQ/cd8ZC)#;EHV__HIe>5U4@+1FY/47-;d_.BHV2ZN82D^VSd
5ZD@Qg(UR<b:HT7>)IKf<HK-^FR)ZfF#HW,<=.:M6ePM6>If2A7VdIeX(>bcARB/
OR2Nd=[YK1KdW,T#R#U@Sf>L//G]8UZRdH<,Q04,9-OcQARcX[2(M/>4LNL^K#WM
T6A@be6SC4++9PDLB5GE9.X-P[ME_dG-;2f,eO/P)L=7<BZ)WHbVgB8aXF\e/K7c
efFUGGeGe&bD_Ie(/GY:K=/W(Y5LdT?6Z^D7)AP/MZV59]\]X,/<L:B8fg8F+UTX
U:-G>Rcc_O\M^(+G8@aWC(M+M/&eZ@B(GZL<;.)52,)HMES=B=9-)R>?:ZL\1c//
O)2;V^ee;9V9VF&dZQFX=@PfHA5VDV#;ICB)[NQ>Z2(Mc[:KXEO1B5gR]>D&HaQZ
>&0-D+>1NMG7104Mc5=g/68Tc#:;1C)T76#AE=>Y5V8&;XKW(_^bg<&6[.KD:XO+
ZAN-BN>+fHH&Q1M/I0EV?(/,OcgAK(5QAB,1L(dBQ6#08#7ddJ+BV.cYLOZM]dLJ
LV<RM/a._6V[^67^>J2)B+M,0d#b9XRHC4BDSMH)92D9TZQNWYNa(bP08eK=&R6^
58Ma#YbW[EQ^=DE-6cATBEOX=YGd<M60IZ1^0SO<6S2gS=f&81(5M:X.,]:M<KP?
Vc#27+\NKOa?fQbOgCV2C&K@IE#G4BF<Xd-VTd11dK<NdDNN0K)Z]HeV^(9dKN<>
HN_TH>2.ACZgCS6+G.SI-1d+7LZ_-)2Dff-a427Pcga(CU,#N(2=RPP^6HF)d^0I
>NRFWCMP;S@f48L9b?6VPIJXdU3-@]_.<NU7gH)]aR)AZ&DX<Uf\R2R4cOW)0C/.
bI@3SWHWXNT&[67d[+X(,18a9a5KB_<787O]Q^1T-[g&]GP9LR9DS9e2WEd.,cgQ
<O+J3aT279F(ReUbTBC,N49NY?@IRUFF=D,g3CI(2KZYJZQJM9Re9SMegOX1SFR/
/LLXZ3D.):cZ+:_]gQWJJcgW&(:P;0(=U:O:C-AN>d,:@H-#@2X1::P<LITUTW09
c.12WBa(/X=8fca7.,Y,YIMOZF)1-+DAS&@<WIcF.T5bAcJX=SJE/7#cE68?E[dE
H2E<cf(=W=VI:GQ+eTZU^1ZZO+AF<C:G#.d=FTY,EE9cUM(\^[;\:655KZ#NXK,b
]fO&SJ1F:1>d&U3fL9Be:^(aIP86>2M&+Cc6(.,IT0UW71JVgX16:9S=B)-0aDF-
GS?+G-S13UVO;@,PPPDYVCJ9X[K)6gXH;)S-MgN9]MSLO5=4UC1+2,dAN1B>78g?
04d.geca#d?2?d?aIC(^KG=]OC9E+R&T)GCDUIMH0cZMY>AUAB.,R-<:[#]WXJa<
Rb;H@)F1&4OR)Pd94ZI5CEbTaBUZ:WBf-;UAGa]].;Zc9_^AC4E,[9L0;;CSJf[-
I7<2M3c0#&>O+I2471M17Q,0]b\)6-O]P#5QR[?c_J7(,C-;^K;X93bI7SX^VagH
X7RL0]e,Zg;Z7GROV9WPM);5#=1D>0\OeZ[0AG:8^^bLP>I6(a2g?dT#I)aZVND1
,::J?RL6#?-@O]60.Y?Z](-eWPE@IUZ5?a?E?M/TF^T_X.<0E,3c(:H[[6bZ-H,5
HIRf3MYN8&.e>D=DG#[U_YSX&=:6a;:3b:VT2Z:OB83E)9Af?GDH<_;_]20@eE9c
[fW+X)XV)G:QWC-4I2=LbNd=&Ca8G:+R7BAg]=S5cO&a^g)(/;IJaV6DN-^[,F+L
c#^<=Y,9UM3WbCDF264V2H/;.XA^b2H[WS5XZ-ZI:=O#2dSV@7F>1ZMKM^B?&\,@
X&:#(B<PRNFbAf0,=Sc1T\TY4/?6[e5)M]4XN?D]T\\e\\K>/_TfBJ;[8gD2H=DE
[XBdVB@TDcNL[UgWQ^CB#XE:V:=,bU1L9]FgN:W+//a9_Z)M#77+AJdUZ.8WYO[2
?&1(2ZAEIa@a0aT.Z0B#K?<_G0A,Ic]5&A0;N??bRPG@,D+:-9<D>IJ_0T+>=>?3
D3Y)+G^fD[_I7>>-eW=[eCU_4?,EIS_9?Ae3L6M^.,KCZZ0M#I@VZb4Oa.JVfD93
9>A9VCUJaNf1MP>OC7DZGPb3H,T7F5M-J948?T.(Y)CB(@R9[&\=a]Y9:bAa8,DQ
/H.>MgX2;)V@dS&,#SLQ)P045YUN^f^G)9NBYTI/O>-4/eaJ)fL\,Eb(;V1YF>&,
.IcGJcM-&^,3aM-^-X>82E+:?IP]_]/6U:dGBN9aF-^f<A;cXS1+UI?NL^?I-Z:=
=4:1bKFcE/B310SP<J9>^cE/4MgX7]FY)L4+b(UfB)LC.OZ0XK81SLP^B^&L78A[
0I+HTVQ3K:e2(CRgO^.8.9IaJ?U9T7U/M8=,/IPXCa?][M2DFVSc8U,TP/=f(VVX
YQbE7(B16A;X4B^^-Y(c9<K=]#_P<c[\^7dC1-3.3CQF#afPLY&;0;J3;,;9[D,.
GM_RPJ2a-g@R.861H3CGUQ>=2b0c@9QPcAU=>21)89+Y#HV_<b_4_N?_T#CaA39B
C@Z>?VfM^6S#CKAW)+Z1/\;Vg8))8]SML8?E2(2bg/HP_KWUc\?UTCa1gL1f+\2]
=0@VJE4DLc^+\AQ@V_3D4TaLP08E/EQ3&Q:S(^O>4Bg2XB)4Hb)MQcMPIPNT]GXP
NKS^XZ:O\Y;>LT0W^)W\2)7W<.7]]ZU?U>D?^BZ68@D\O]#6=aV(cN-@Ac<,5f-Y
fBDT+.0?\GHR7J^\+A4Y#JN@7_()<(UPTg2U9f<_/N<-(HNU.\#)K7/Fd(_VCK_Q
M6B^TCQeT\];cf,3408D:[N[\54&>&b&#:fT0K,-;#bP#5cO=Id^QP>4OOY>eEEb
^Bb[FA)[Xb-P>ZDgMF+ZNW(MRb5)6@Ia:#L0<cB8,fGAfF=NZeX5UM/9)89ON<+0
/Z&Je7UKPA^F@.(W7g;=^.4fWDW:WgB]6fEb04?@1F+-V:aL.-3T-^[HA>);c/E?
fBJ\d^(TT?(1,d##=eDI2LR)5d<+N&a7_c2f:e@ZbW402I0]=0II0?A8:>d(Q7Y1
ING(+QB?J[[XgdaQ&1-3#VOGU\6EK2_Y#W(D1:+=)0XF:\Bc1-/0O[4>Hf/M[_#Y
2J5)I[bHR<?YQ=4.)8PVcH&K=V3A-aWFJ_3YIF7XM2NV9F/)+W8N(JSg==\HNMD0
#BV[VHN[83\XTN=P+g<=H0QI#d,F,Q9JYU:.NXe:65:U5POTH?(P0.ac\6A)Tf1Q
b@+34^U:3V2^=g]@3R+JZcWL]W:E9+f_H@PXePdbX:K-ga=_>RS[:P=+Pg2HK[HZ
:##aS<JA#d?G=5\J3GLKSc6;;R:<MU<SGO@-4aX;^V8f6QMR&IK<<H;=.2O4:L4.
>2QHWESK988@AVa>?BIZgebR4@1(=^H#e4.;-TR.d^#];1RI:.Fe[O?]QG[W@C6;
84LMe-BF)d8J+4&S.NMGBX_K@-?]^Jb>?dO/LRN3TE7RB&Z,+1LCDOEf#1/I>AG?
81(,7.,ZdIKF-Q:4])d6G[QWJTJJ1-?R_;\ZUc[V\C#VgK]X-e2_3B+gXdC?_6dG
D/:;N?.PHT@f)T.c.HYB1ADd&R]Jg.?O?(^:;A7RX7&^EBBW0Qd(W;7NPAB5WS0O
)fHJ^L<GTF<B;<6Y6)@.&^/.Nf/eV^3U]E8A1()a,Y#@C4If#1:XE7>)b#>1.ZL:
6bC147M+E9CU>e?da95f(cYEY+\[EP&XWN(QFY>/Ff80;e-6\5L8g2RX7g0V([Mg
H<eBeN^S[B:4US0O)E)3e;SO\][eeHg&c=&#A)[8OC7S/a/f+G5WaE(e[A>@7fUZ
N9S)IF=2BdN,7G?0]<=A4>d+ZJB+DSM]f>G.Zf(+9)IcD,fV0:X7EdS6>09IM#C0
f#bgZ/g5gZe[1ZcJ?fb5,?T\e@-F?#c+YIJIZ=cY/2:2W:dKCG[NVVDL32&RFY6e
-(-,6JIH5IgcY/f0Y1-\__[U[J98V@^cBB&5IAQ<A)LVUQa.^-DDPJ7F+6\2A.6G
6GL?.09b4_)96X4D1)Y+&V2fPUT=ZPd/L4>7[_CKb+HSNd^G#OLOS:[T0C_XP_,L
6PZ6&R>aKC^IfEDRG1.gH)PF=1f+(]L72D;#bSR.RQ+D5(TBc4&5JQ>O_b9:.<Y_
:8_?>MEK05g:?aZ\c1KebEYB9:;?;MZC@2KA&W,a.@Qc-[[/O\YT&=GFABJ;H@g>
dQM;#_=>B<cEfL=)6SWL#NCd5SNIM(12???O]?4M_LFMb.EUD(XE=UUYNH(?4RF<
>8OU0Xg_6[UNg@U+W\\6^K^>?LeOTe4.O?K-2.Hdde-.GUNNOUe^K1L(MX?#,N>d
PUVF5BAbF9TY;3LOb&)VT4ROW/Sc.TDP[MC.V)KWS>.5_)D@()NcBHWF7T[RDZ/6
USD](D5=XG&]cfK82M#9+KWEEV6)1I.<MVE7#_fO;5=0,>b,^c?C&N:BVTIVAFM0
TJRbNEbS:D/1ff2:B062Z#O/I\B9CfD7@K-:^#e/Of&PPSWH(fOeeW\;,1FSZ<@;
DIDbIQC9OR6M+2ZA]ORe#_f)>;/)d#J\g_eE#VC_TdC.ST>(TMBN^Sg&?I2E7C#^
HJ<7KX@ee>@@X9ZV-D[PE=,-XCS164T:;KSAGg\),Z9_@,e=7NI(/MB+<?&5:#H-
43Na3WKYP0N<cd>&K;JLdO-.JU)e29G8>e@L_0OJ9V9]gNVXQ:[/K>3JY/A5R0&L
6&.-^P&-)I5^cZbW4]Fd5),g?S1eI0Y?5XNa8d?ec_<Ze]DF?@d\^2a,ZMQ8I<?X
c>-,7,4FWY0@c=5KQ3CgHQc^Q&JNP@fE_4fR4Ka5f<ADYAc]:J3+WXJZ3J/EV<5/
DN\6f+C38Sd>7A/BY;80&AL/8,3]bAI\6[L[g+#/e>RMPYK[&NDTZ?XaO/XY(>WF
51:ITYd(ZWaZXW2U^2F5WUb&5<3.4F?;LW)3U16X[1W:6&g=L.g#O[CB5O;&f#US
(GU4-XFW/^P5Z9@;:dT\]IZZ(aK.e-U]>QadbN4E#NOcIPdUD^;&HMRA+3G;^(VD
efD&@?.=GfeTYgIPO;>;&F)K7cO[X6faX&7Ud):;>42AaU\ZaD39g?D:(\fL<8f6
H.BbW@-MXB=(Fe4DdS@fd]]ES,_/C=XCWDZ4g_0XDAPGW3eVX(fE4fQWA)VTb(_X
.N=X266RIgLHag8FGIe+NN4)bMG;_GDYCCYX-6CD&7/Ha,2d,VA/<fF#OX1?FcK3
\M-cYJMHfM.aD[9FeJdE3_ge9bLK/-CPD6?cQ^P^2Y9<U[4:<;=0\I]OQ;&>HE&,
;/:(B\1]G6b\&;F]N[Zbc1PR;@Ie)+MdaP;/CRa0>D3J05>9P\]L6<QZe-@IHOMR
dF+\>Y&7e38gYQ8W-T&Fg7TV3-V7d;SdY+=?Nc&Fd1Na8-,cE88#WBB[Jf^GeHBV
32KUDCA>2XdN,,R_e40&McQQV\Q[SUee4VO0eD=&aKL46.<ZZMd)K4QZ46I+e.HF
97S9:@G7g3U[N8?)e\N?]f1-XA[@,@0Q<+]/TN9_JQZ:;ADcQg:9,;0LCP^E3O#Z
P@Q_HaKQAb</TD[Z?W[0=HH_<4Gb0N90BHO51Nd^F-[>1g<-93TVcXe-<AILW&+I
6GTE.,MQND9)6JVIF]@W(Q39G(bW:;cQ\:fLWQ@2?-8[\^#:_OF(R0TT&#PZb5Q\
J?G7\Y1#UK=X].+[#JPfN[#6Lb6f)+fY3MOU9\]gM?+&&1F\R[aU04=EB^DBNCD,
X)2QZKf47g.?_O=@\@]RB7B->3d<g<@[;Q/A4E1E/DaTU2YRUR>@=5Ne2?9&0fIE
c=]:NXEJ4a0e6[@=<9I5E.4@VMFa0Sd,H[J5_>>@d:9O92W2K.eWRQE1(G/#;gMg
adeFHQ<Q]L-]D;bND9Kf\GfKN(&6:>SS;7##?3W)&723Q]MHOP#33d/<Y1JEaY[=
P:eEGE?#CTfda)b1+\/;K=12(3B#NFL_(7?eZ[RX:H6d;aZbJTRW-<c;/WD+e6]B
H(]+HeA7-_?J#O4cAL60?1c,Z&4cea1]#;PT?-Tae7>G2C@1;QgVbTPAVZN5Ef]c
gYT[A_UCe06=G<R#54Lc[45aNZSQM_H8/B@IFcEdIe/eDNC7N?dU?6PB77eVL0[6
9D.8;1>fe^OTG,35cU[H>2bA_?[WU)JG2@W&c#K,#D;UZ&,TU^Sc8[X^Pf3;L3NO
KPL)W#:/N::8Q8>=,CW&YD6:5KVR5a<:6F7Gf<b;6[)/Wd>_)/XPC(8YU5+(c;0Y
Gd=1]T6Q+CF7FW.YWHbO19<^K\M[>XWR-^\FCPIKCM\dbV?:X66&NYNF@RT8AD_+
#IV7@aCO\6&=61>_ScVcfU1XD@Q-[/K6=W35&6_3RFd]MAG)4J7C6L0b54.@(88@
I//-Ua5K=@<B1,MbN?7O^1fc3W<32TJB:eABaQDPDOX856WGJ4W_aS68ZHFJ<Y\B
R.L3EF-;DKQ[Z(-Ia&ALH-eV6B>T_)=Tb51@Q1FV;=JQ<Of)+g.Z5SS+WQ1/69ef
/5YI\/-d.)<&2#9e-H_TC)=YZ[8P@3H3W<NBP7C7DaQ._0P=dU=)AMQEa3Cf2_<I
V;P#(\<#+/(\HZeJA>SMNW+>RaHP]Z7?WS?3gR9a6_X,SC7&52.E)U:NHN4&)fY1
V..I1;[V0:dDc.W(\<&YVRSJ2OFd>8\[Z,^3TT.(5K/9(]L(?5/XQY29MX9KV;,<
NWJ>G7NXNX5+,8=I^<]76CZ>gZ+B+^8/7YR+A<:b^.\GJQX)A:Y]C^UVKg:K@UH.
QKV;#Y@>Z+-c@3g3M2G8_2M]WV8XJ;R.c:f2T2c5?=T#;YUa0(Y2Q=[e=SP[B^G)
]H+WBIfF56NWR,D>?4WK4V9[aIXMDG^&[-3f<SS-))cZ&BOE<d]Nb]D7&#5F<@#C
8QMCY7=#L+gaW;C,&6GKNV_38UI#N6R5GKV48^)Y#@K3A=ZA5K>3:f;@TG\&2K[]
=HQ?\W>-25[WH8-/4,=R?.e>F8O95.4=U7.M+c5HfB<@3C&G)\SH__8R=OL9SbI.
(>a6]U>6\GP8-FO[6[=TT43C8LS]U?4O?3EIM=FBQOdeVG[f?C:7SW4cOcF<3WH.
@FBL19+&Q6g=EDa@#=_4_@RPC71VF5ZR)Q)@CSd+ML5IAPOYf+Kceag84&ILc^1(
fFQ<3UDN\AY@7CIMc)H=MQ1+eRPNSbd9K8eGKafRLdQB-@]DR12c<Ofc5QUSF96F
K1C_>D0C>LJEc\3XN>YW?/c<<de)bFM;:b>+=PM9RTZ>bWWa8O(^dUb2K,D][5eQ
5?M)-.7U#UM<Y3A3aU>;/RE)G,PU<L@&@=5gX[00CWD1LV:]S7V.E\beB]<;NUX^
30OG\bYQ.(VNDA-&2=DYC6,K6bO-CL\H2[GMAaU.N)D,Ja62H)44_BV(Q7KddM@/
&LGbE7DbEK\/Ld5))@fK6+c,53?W\CPLO5T[G>d2c[D[99#AJ_fd3@0);Vf+3)RQ
cXDFTH@SQE&5E>fU;)]9g=,Y@\1K&,QeAWS&Hf+::^+P=cE]F=LV/<Q5a(QP(T5a
VEa/@Q(A/;HdG)NQ(01WVfR5Wg@HWB-9=YTCdW12&63+cd,@Y,JU&1@#EW@>=W9M
)7Z0H3^a+@06a9[GM1^)81(?f=ATFX+a+<MHY(#I.@Be5P_/>Vg)+T7gW67T<2&M
#@b8V3D<:0B0PM;X66J6HX?S]JP_f.),Fc:@FY>;4-;B7f@=H:I4W=QR6Mc@QZO;
-#Bea].^9eZR>6f,A56(G+C]P(eYHg_R)<<Xe]BP6E)V@]QNR)(LLWTbU1HYM?85
.R:JN3Y-?T>@71(-&>4aYSWgDDY?4K=)R]9GCcZ7X<#.<G1VY5+J5D3&AE20JA[B
YI[bKcYL;?\c^NH^ZS;<g4EK7]T5XT2QB8<\g\Gd]+86CVTMKQcQ+^a5S]ONbKN?
=a2<QV4,5/9OKTR2-<&>,.?=T/N&8&Cf=-cUd4V2<ZDH>f34Ia(<Ye(;JJEA@gQc
Ee<RY<V0B35.@_^<f/ATWT4AE[JJ[G&11X7M,@9)8<3QTK)Ee)A8T[#1&HAa\AM4
CB:TdBX5DP-.Y40Fc\S=8^=4>Ca:#7-Q.5^RKFb60V8Z(3[\6L,dHHB7gf,3,B9^
=5F)#9LOWWd8e7-.H]A1\K>J<0>Q&K(X8GV9F+79aeRSA,F86/bP.@QR--E[Bd^3
KL47VgX)>04W4;-=2&c=RY0I7d>L=V\X_0>=U7cG4VYc5N0@XF;cUOPg<=-a8P<8
Lb-U/b=I^L18L9]CaQB^WH8V1/4VG8<KY5+9<R.<TN&dAaR(:XU4D44fO@9O^9N5
GR;+[J]=g_A)P2CaC1X3;AGW6]//XW?YWQWc1=W]Q__DcGeP2@NN3Z<G2Ja)TKUg
A:g:bJZ+a]J2D;L=AP+<d_fN/EDd(D/X4_R6dOVfTFZG87Q[-<TOL()UTb^c?T+f
g(ZUJ0WV+]#7[dd[FN@b)8MYU@\8^PA#164DOSb#P>CCR@5)-b;DI:.I#8g2J8eZ
&9;6=JMMYY_e24(M<()G?L.7OS;WXZQ5fX1(#=)H?6fSc9VGD-VTS3+1]_ZOf^YE
-]ddeF@25_,.9YA,472VF-0c,CP3a0A//>+X8N:T&5eA4gg).-2Wed[5D-#8..<S
<W5S\/28(6-OKf?IG6XL;c[,\)eIAZ6=>RgD=D8GANO40ae#NZ9P^;fV//)NXA+P
UJ5N0A;M8\K?cJ50EGNTA#^c>[e=G/C#<cJYaA^/>(&8XSYcVWa:Z94H?@SIW>7R
UFac#58dPgD50Y5VG;49#H7eJIC^[Md8a5g3^[]7,R]OL@644JV9O#FdbcAAJLN6
.XX4V2fZbQ_T(:MbZKR]<=[1>;CH1N1[NcC6AFR-[R9/P_233J06)<YX9c),#^N+
+,aeRN:2@C8+266COHM3bVPC5aB;e@=Q:6.+X\TP,Mfb3UGg161)J8>a&6aO620a
(@J101e1M))\EL(HU/M-#XKD.>Q7W[8YT]CcTaI[\N?)>JcgC.e]X4La3X7g\6^g
7^OMIYKOdK,LZO^bJ2.=#K;V?[WVT[RSKF;.NL7PDHKET1T1dP[\8J7E]VHKR0GF
IUSd73;3^D7B7KRKP3):\A]e4X.@5A\U4=HeM)ARUO<X&7?#Zba2(2L3AcZ)@9@3
N0Z6/gYLIE/eW:2B8R7eKUW&a<-,8e@HJQR;(-SF<RY,_V0AKZ#&H:^D(,-9:SB-
Sc]N-#02=8N5MO@L63PBE.P:L4SU.K2.&bY7@)L]/G>?6U@#/BeJf?E<H)=g=G+?
;&?a.&bB.MI1CD9.M5:R-QA2F+gdOQ5G(4NAT8;+=B#,gIN>C5TJV4,0L>T8<M/^
677^F3G2-Ha\I,[?dcd4OfCR-bK(CCa4N9;IT7CKd2S/NaR7&4.=UM6<5EM<:2B1
Y1.bTBKAK?TJGSg+fOPT^\&_5Y=+K/cRTegTgM068J?=+FRBeP\+f]aG,EgVWL1B
Kc8C@NEg@>02ZZ+Mb;G_W;N01P?JFg/df.9?XEUe\Oe&.CZcQ=O6HcQEV1b2O95&
Bb@fL3d<IW)3)SP>]U/_Y_HFB17g1?=/6GRK8>b)O)PQ5\)6/679Y?P&OH^Vae)a
eZBC_fX#b9L\)V5Q(TX7S&Z8FD[G)NW=^A@5dZ9P?c^)>=6BH+VcPCR/@+C+43U]
8;H:ZL8/PWWK+36NZ#.NE>(K:3&VE5NNWd.T_2QX4-fVSCGeg#Ca]+B<70CfV;I1
4NB<2VI>aB.X(FUc[N>F4)^@gFU5@W6<^H+?BR0X9+7AH?g9IH1O]VS4R,8XPIbJ
E;HS8]GfeQ]_DLgSDB?:KQSDC?HUO(D/-U)\]=+#,.#T67L@YNDEE@WN3UfZWTNI
X+#8>7B;)&4@DO&(0(NUE2P(<_IHB<MX5:WA_KY3O-c0d+U5R^,X>Nb3]+PHQ&Eg
L+:]^Z0a;C\4SH06SO?[]IN.eEM6cg7?F8I_Pb)WCaKP_\N\5DH9&^4T4@UM8EZ]
C_DAJH=QRS([141U)I\5\ML\#E-f_6b):;B</W+[Ed7?,G,Q6ULC^F<#]d7a:9UO
&S<2B<FLTa?[(;eAKFRU19QUGD50[@C0eZ3KK<W(>.HVT=\#-)+&,@).[a5B@/1=
0D.,:Z&&HMV.JXALP)XK(afJCK3a=H=KQPM+(D?NIf[&^)(:c4E8W4)BgE<IOLN+
GbER>JU5&4g8;APY-S&M0U=4D)[b-)<HV0g;04WI;_AR#a:0YefH5LK.?U8(<+c7
[6=4I[K[FSJPAGFZd#CELU1M&EVZT4)_W.e8=7Jfa7CP0Q]->d-:&aL/OE3XN1_T
.3_8I<YE(V.VV\QPW76dDXa65/YSPf-[T.<J7YaA=21U6XHP;JOQ:6\KbB9[ddBQ
Na8aad+gYKE2DA=9NB1dYI)EK6g-YTMI>YCFOG_7SA#??GI5M=+c=BaM3g2fK#N&
/QW0g?)#@f5ZH4(2DXQ)[\HNf3RT>19WEGCEcL([gH?IXXANT2(RB-0VOdSAC-\O
17[EGe)<EMd5L]#^=2)/8e5ZGXd#:HEe(5<Y<EHEd3V0JDQLS#03136>:V>)6SMa
1UBG:NE=4T517]3?3)Q_DIU?9H79Z4SEPH^KJYdPZ>,<-?0[\GF.<:4.X8d7;c<R
HFUFB4P5#9DbJR#WN:Y3HXN<cA8-.9(;4/FLIc:>LN:]X:4be@X0aSZ3@BZD@e2+
&A)>JF.+8@\))cf8UJO=0DE4Sbf25Z638-PfgIHZ]ZZ?9HFg_TCOWYe^(GL378PB
ZEEbPWDdU<CCCeA9](9NMFR^b::9;^[(O..8HZ]RB7a),;X\B:DgKWcMC6:-:Bf2
SdM6+fb:N.SE>0e5)/[P^9.5FK?R&)<)HQI._0DRK&?H8VB35Z:7O3W=<7N@[TQ(
=0)fOcQHES\RX]fdFR,)[gR9<)2XR8a_JB&X1c(d33(&#/LHNT&-C=04MUQPMT#b
L86=C8OcZ7Re_5NQJ6Vg1J/W3:b2G6F,D_UX:5E&UGDAZf+++g96DT2fG0NG=05X
KDNX+#L=H<WSQb^G17:NbESRV@a/LL,bQb(ME9e<FYbA;<Ka3(B,eF-LK.01fEPP
8eLa[:aE3H7cKDQ^&6ZFcZA:Y<1e:2d1,Hf:S-Y3-U\9XATUG\De7DKR@9H_DG,.
+7PLF&^>6>f.XHC;=cGE1>:#2g\2/V7bKg4QLGaK>IP9/3_/EOL28S2XW1:<b-,/
^_3QCR-WI7dU=,-Q)^K\+N-eJ?g\M;aHfO7N5#S6aI(@H[5dH8F?=O<#?:N#-fK9
G7#8dUJAYa(d3MN#\+_>-QE=R>RHX&(#N,L(1W2X3>^3X=8W@95fa\)QRB>G-f_-
L=2/Z1B:REQ/812fMRcZLT9cO.eE?[<-W[=G[V2FPg+RWVO#)<<^T0[<VTN,_QL1
E/GOdgbG+:[X/OIOKXa:Qag+N&#]U.G^>W;K2>.P,H(R@[-.B\-+-ReY/VIHdb;R
>,RP_U;F1,a6NFQEV1X5SQ]P4[/7COWOag<dG8?7[>\IVgX@8Y5G&Z?\UTaD)bS6
#U8:OA8LN[AOXeEBEMdc3>]5\TcI3McdI@3CDNNf]D2<Z9=E\<QR8+R.#5WMB[ZY
JE_/7&\YBbB;+Ga6eJRgaZO[.X)48VN>#;5G5A:VF@+XNE5(N.GNTLZXZ5&HN7]<
)eD8WHYYec&QUAgUaA5[H<A6+FV1f<<[dY64+NGDC6Yc1K\)+c.6VWV4PXXK,g<R
N(E31VDU^UcZ:gJ7;G52/IAfK/&^gY=L1T;VW)I5^@/+\QVdV2;Xf&O1Y&_R/UE2
O:c\\6?U#5YSIL@9/ddB2B+9\Jb18001BV@.0<@TK#]>9),V/D[>55X]^L,c0W)Y
#:FEa+A&C1GGUcP-++.=/SNQT/G^JWfM+3;;.4PE(+798@GV-dC1MXVSXJD(GWS(
<Y7H);)@IE53;]F,WfSBZ2?F\&T9ffJ=b+1Y1Xd#@(Qf#>.[0HB>JJ)JI^9<>[3a
S,aKg+=T3?VJd4HUaNZ>D2.<U_7cf\SM\Vcc6\,QC3:6(@=fF[5dO/fXPW3RJOT+
9B_K1279SXN3#F;fYHO#LXdB<QB?=U_V#3@bS3Z4_2SJA43(Q(Z8(6UN<EU=H#a-
U7-&5EW:<Y7JZW\e5YH[N/4,bHC#a>O8FX\MVMf:-I4GJ1/J3Lb-#5/U-3W_0Wfe
NG8?4T-b&dXC^5R1S9@b7(.c@)+=[K(/#fJdHW7DB]YN&ZVFDW8Ce;>U]Y&e7RP@
LI=F>B5]R7gMWEWHM[QCF2N/_Q85<]A(K;@MJM;\L<=7_d4g2eCLOTaeHY08\eBH
?J0=9e@6EUNYL11M4b:L35:OJcP<fa-@a5GLR)8,#DQXZ=-CAWS3[Xg:4M/)]5RV
8?NfEf^-Q;-[bfP1>2CCQX\E:Z5)GE/@NR@6<6Qf?W)d4.NFZ3NG&BJ-K;R9Hd1B
SD4?>KS3A&,M^g;SF,-;KH)[T_D6G3S:eFOVJYY82Q&CedIP?9EL2\XB&g&/HD[Y
5]3WU&D/Ye1EI##ND1/-0#@0U[_ee4)-NS@BEBW=#db)P^)+0[Ne86QUWgVTbK+#
a=<NYSYE@G^G++ZA&WKgY[gS8?O)S-U.L(eZ9CCIC[>b(]F+[COMYTJPd>cSRS/K
S8D,=_RGS<TIa^H,MU-bW>T;ZN9U8E=5A-c)EN0IB_TaC86NcCLL2eM#-bWR0EH=
Gc,PBa1cYDAUZ;U9A^Lc-W>b,AEC)H<g\UP_VeB,DZ==^+e,1@2J>C@:W;)^eF0W
E--T-BP.M5NEIL,2eJ?cYW2gDGJEIPg&>KFN+>5<A2QAZ&P2IO4?9F91<<4JE(P:
[#>KTU2&f&:XEY-Ld6a1=9f1>bfYfaaVI,3f/&aDa\8cSQUS^=E]<0M<TQT>fGa\
\G4L.ZI8E=SO(BI^Z28_.>6_T<PPX9-3#4&418CE);<4/Q<]Gf,@=ZFA,aX>4OV>
C@\X04J&X2GJJOR>DN.E4U#2,Pb07dLLQM?63=2^;JNV&UM(34K;)K.?;,Q1L-^+
0]BJaC;1\7<PT<>27#05Rg&3e5eb]V)-CXb+9_;O7+2,^,RESN_2QB2TJ^WUB7+W
R\f/TS,Ga=4U@bb[1S1=2H)NY:?\&GKe_&c.GT<F3eU=?1;UJ5LNT<C.4690O#>J
0MJJ[8R[0/JRXDOEA<M[K5b.-Z6)&(19FE_#+RYH2KWZX)?L-Ld57,7Q7,QWA8?9
cYOGe:XEdYN]XVfL6c:MY/1SI_UU^MZHLg9Y_MTb^.a:>(L;)1c<MW^I/7f4&2#X
=c)0.A^/<LY7G_FSD(V9?;cb),1FN[E5YW:S4W)PQ@5I)F_GR]6-X_PLSg[RAAG)
5EG?:UdX-A(I;+Z@NV7UYC>b:ZX2(V65G?PSdaT^]R]OIT0CT;aC/:<.+PgHFZLb
K&63W_2-d#3_9I?G[+J1I(>Uca@=F2O;U<S/K+^U+A<g9R8.#I_V5EJG<I631b3:
FZcY1-\+YQ<]EUN,&R0O)QQ33QVcNZ@cS\J8PTKK&UaTI).A7A?NQeTKS29;D;U0
SWCL\2_N)b7@1C36+6ES&WZJ5WB=+c@E0B@?U&d^FXbLcO/>(;4@\^1FW@RXOUJc
fcPIE:QdHR68BICf+_P1cbKU_##IOW7-\S12;-<Q@CY(8[#L>(CRb?QcU>T56O(]
4LJSK4d9K0_1(#Y_F8e^_WE0,O61N0SW-AeCFESR@MHfQ&<S?g(6/=bWgc<62(S-
4b4-ab.]V5JeKKNQ<0^403@J?]M>b9IZA_eNP\^AIC;H(F:9SRN)X](_9]/G4E#:
G,4<EVRD#g7?75c)L]:?V<55L6(d[eV\2\KFD?KD@<Xd<Z=T>-H]5df&+=2aB4=;
^aX4)Z\K0/:-0&T#O3BgXAWfM=,D>R71-)IQ#>CBC<?KY7aa^V9ZeWgc-a.JKGf,
3Z0?\V=_/SLC1ZEO6W3VQ(5K\QS1G&/?f>8g@VTKRX><@bTZb)P;N9YO7O<=L\:-
Ze/GfXRDODNW<24e/<^T6A4UT_XTFdCQ[L5O:gM:3<9NQLEf<N-R#gKJ?PeQ6H<_
2O-O-TgKXg+9(-SYg<0X&0faQ]&&BB\SC_KC4b3g-?LZAN/67da-ZBJCf+;SR^&>
-[_/R-P9T;[FDbF[PB0T^^B/P(GYDJO[E?:7+1J::ADQYQ^1>^Kddc]^X0F,bBBg
7MI?=Y)>7b9IVN08KPBc5I2_#_?f::XZc]WH&A;,YLdJaL^/-XD9VZG?+6WgFcQO
F./IQaQFVXC>\7:DXUICI.TSO<EDMKU(JQHVdDS(VN(db,RC7^2gQ\3QV4:U:XeB
be.TPUR#c3O#NbHY0Q62Z[@BXPfL,8.cIfXIOb[##P5+8=M,<Fa/7-;<(d:Q8HI)
0)_M[O8)O:3?71&D>DPZ<AU9b+K8[cY]]11NcQU\H@V<+&<NX7L0c_HV5+:/_P1Z
,4E-0KdKQS;f5fBKI+\-La/^CJSRL4J:W:I)\cMJ6H0]fI:H,31I)D_?G5;>FI(X
N:+g+=/F3R]ZTNB-^:82AaaPYFcJ\288?Y,])fUJddORNCMZeUa_B5;a5VG8=agA
G-Lddc^5)E.PV]A]Aa4eWRU\#41UU_bA#UJgFAK.Zc:ZAL<?>7_#]4YE702A&HdZ
L)ZQ<0;S8e[:1LQZQJX]2d:II4M6=M-\HJ^T9K[4QgB]:IUdE3SD4SF<TF#:QY-#
50F1>:,7&?5TY^f^ef1AL(#V]H-ZNFP2JdRJ<9D41#D/3(30AU\_Z5/]Hg^]P--[
a>T9VLODC0GPJ,Nf,=E?Md:WSfE\6;^A,X;5B+8.a2;2.B0)R&5X4=<=JN(gULEe
0^dL2LS83f52>W)=7N4^SNMee-\A_^geXOX)I9@G1?GM;#A)(g-<;?<P+/0;9e]J
:V-0U8G39RTd^Q99Cc4W<PV?LGFd=6Pf2L(.g+<1\B4U:?:7N8UJH([TdO8=ZUI&
5/d_=e4X_>5=JC=T[(ZD/7]/d[BSLB#7fBBg^3?J<T:H8?H+_La5P,2Ed#YNa5F2
Rf3R(c(KY#_X9Q_1M4bg0Z>:\S[cFYfb<7RXV5FQd;,;BGM\#^eBID(Z^Q4RAI?B
T))<K/4[,0YNS.RVH#AD:Y-T>50fbcAGUT=7W0bI<7YRC8M(=#BMUKR?H)=YTT<Z
Xd1Y6a<G1:NFaFTFP1)bXaHEN<;:_(>-:JLeedD\PB]\KW^U5?7gLXA4J06JL+/C
DWAI+=D1GfeX^6Lf^KV_YHcZ;1N+Oad(d519RHeF3eZWR&aCNaF0-T-=B7e]A9dG
IN>1K)SXgV8I,&M3BQ5(CD,CRDJag@EeTX2]>I2<ZK>2\P.@YLCLQb<b-0Gf4#b1
U1NaGKP=+9eSTKB^CO6J79aeW;]<+)K&gf?,SCVa_L8R4Ue\^WbgKZXH:7N01b;9
A&>cW[2f<<K=BPZb/<:8SX6V+MGf6_]OT#DDaVSTDG2RHdYH+NAe3(,O^G@SUU-C
dT,)O8_d,?X4dR.)FIPJ&SC^+(\(IOG@fQ+X/+_F9<RS9F\]45^c#7<(WZ-<Bd^8
[=?(,NYPML7g^P?X<6OL:>U9Md7?GDR[0bb3-[+1TdYJdIbEAQ;T[^][)LG6+>1Q
9I++eNDBR@FGYY+YZ/bceF7]Y0-8;>X\c)@\c5c.f[C<BH#5X,<[a&RV@H)6A?VC
KEHO+GdZfc-)J;X<GOgM@S]VBX47/WdH:BfHM:]S_&QTV.K=L=&/ERK_Yg>P:).<
#^BGB,9FXa;[^N8?7bU#8,+1\-6ROI04V1W\7/L@bRCWEPB<Q4S7cC@b:Cc2GFZJ
ZLeN=?^a)D8Wg>TB8X27N^SL1^W7.g(0[g0NW#dU>9]YN2+b1[C5&LI7\17E[>_L
Cg;^CZa),ZV;f@^O]SWH\3>CPaa-4?+RHW\8KQF=(;cU(.((-&-/AQVP:a+2#H29
PE+T8EG\-]8IBE914I+BNSJ=M/cXJ--L,0?>Q;a0=L?NcYEGW7+@<@F=\;<BSgb6
=87<S^aH2+)8GV:.+[&YRB5GU<5_1K@;AT_ge@4g5DY]S8=[YD,aRD6GZF;(fa?e
PNQ>&4@d8=@E<Ma)9N.72>1WKV#51E6LX)+]d)?EU8[_C&dBcBY70DN#.\E;K9_4
7MeQ?,VNN;0<gLf[U-1X2[TZcZ+.&[IC:c^+X6F##_X(c0YaOGcO[9J=GS:B9&]<
U_4#&ESg_AE98Id>8LNM-9C+e/GY7:.[W)<@(e@@)P)Q9c<)g^gD)\^/</:BE:JW
c_cQ^(I]JSLe,SA\Ub=5Y&HF/24Z>N.SBe],68P69VVKdG;ceg26=LKNffQV-S0C
B8L.UL6^Z\]\8:PL)N-?]6Dg2H1_#QC0>fAG^DTUQWL+0^,I38,f>9L3We/d)W_6
_O\A)5e>9<&VNDb]=8S=OY<38?)&4&U>.g2==X<0ed+]R>;We#_1AT]@e3BK#Ob9
S-N>PZL9[AaMc1#D;IfZ>#dK)A_O:4851_e/cLIa=>/5FN<_AG8/].R>ZbAQ0J:\
>e^P5a7GX=A#=cO/gN:?_6.5J<PX<(&=R.K^He3SO0LF\:(U<KZ4?H&5I54Z5+A=
b1[8&Y7JM10N#_RPX1M36cKAg6P=W50C#[ZS>[5V=C-fc#EJ+Q^Z.^H)=#HeM8bV
(a9OO4@[P/H:de?W1]=92K^[(D9(,,aTO7:MSC]OB@aO0DG0L\O9#:R9SE7X/LE0
(KD2ffXC<LKCfN/f8<bD^dg]+04aC=MK@@#?)3)MJW_8N2AI(S^17H.H(SWe_eV=
PP+:SJg9Wf&)Nb/HdcJ/V<[)5QBYL7S>CR_d0D/fY-b4g)9R@Q1O<U)e49J(31N8
KQcWE?^b2dAN9QUdP(SYg9XP5.V?0(.#(::=8?f\^V(VZffNU52:7/7f.);PQIbX
HZ.27f@XA_gg-)4G,ZMd-;]C^IP(99J+Ne>M4e+<[7deD9WD,,D[\T)@+1.:gHdR
GQCN8?)M.0LY-EQF:3G.<Yb[1LU),#<TBGD0]@1.\R(U>+<Y,)U]U?Z:T?@G^(<J
+(Q2_?7L(X,K57fD@,1R/<)\fKAAKE/59\,Y,147U&(#AQ_L5+ff4E;QL?T99,:1
6=3R^5&1g-IE/^DXAa\3>82X[d?1Ed:#GQA(W?E9a<g#E7<a^KXb_=gZHTJ6F3\(
)>CF?.C&Oe6Ed@Q^Dg+d;,HH6dXdeMSed?FKR2;KbT^7<)Y3>)6a;H9,]\UPK7@-
fL3H&]CRbHcU)bg<\A4D#KQVOcUdT]fJA=QC:2A9b)4S,\C>.bP8e<Z4429-F_?+
MGBe0<Eb+](&c:^46Q=+@<C[bgEJ]O@T+[N&CB;P(U<ed,FJc).<I&[fEKTPgVC/
/(bMIA^P/Q+8f/e@<ULH>8VQQg=IM9-6(X3-5DP9VN9R43+N<Z<H7cNSICgI,?:V
gd7&A-5O?:BHD7-eEb[I6MI],UU6M8,VX79G=<O6.7-deOO.X5IDAa\1Tc(1E0?C
UZA+#X&Z^S@?,/+GeG#C[VP:UP(bHRabG&JZ+GJcRF.=I[T16#M2IOP<M:A)eDN<
_#8I;Kac[FP).K2#D::@I8?@-CTK^^(dUCAN86URQX69CUJ^0;F?<UgRBb?ZDCA2
#MUZ1=cHc:6A88CY0Qe4D68Rb>g<>gf?ed+K7M0#2g[,B5+I/]g]dL46YQ/>[8OK
;@d^U6+F3b,2S=L;.ND//d.:<G+7J>f[N-#2P4R+aIaUaXGg8\KcF@A/B?L6,R;&
f//,a7Ia>>/cUX]LYC6WW@N+)2688ZSeBH5(HScLF:dD;Z.R3B=7Z77)eC^3G]2,
B)>NO9;#Lb]H08<a-[+(IZ9,egU(+<<U/eKCeZ6dUbMN^?+(2I++<gDEA@5]0[RS
;O?Tf&9S?-C:f[NF0CF4VQ8D)+^5Z9M^L+?+XKSeedZ@X7._^,>Ug;aAZRDN&T-]
#X)(PF_KS\FfV)>ILTfBgSGU/-VLa#3=J(OP7<LX#<HGD@)+/)1GS##QKG33&DMH
,R[91UUW2HF&XY)=B#@N:XVgA?KH^&L\59b91TW/d.Z:>L7U071OY4e<<B4+Df-f
73FUg^bY+CeA=PQ^IK4O-NEfaW(9:<@]9?If)2QPMHS<[W-91ZE;Y#5J(@K8.X65
LZ6F2O./V_.VY50\X]@JEM(\?5IXWA\U[eFI,X;OYU7F9H9d,/c);(RfD@7,I&3,
_2D7Fe6<QCMO,6/g8)_>2f?7W#73g<<\BM[?K-/_(8<21bWDgN<;JeCA>bSFEeFC
B<(f;Q6;Ce_YOSNS4PTK8&&4:K;(1,g;BJ,58c]6E3T/0YEHFMJB^Fa/bA1cK5;(
Y1/#MD5/:3KDG;XE3.<8-N_@S(eb(:8L+;6]ZE=^BfB=&g9cOeZP2b(AWOBC;a&,
fJ?ZT1N,LCE.Y_edO\^1,?A)Sd3,;(8YQ[0XARINLDgHce-2]3J<d4\IK(0F,)>=
SVEf)3)B#>I@>&>ZP[)FX2^L(PVd9@E:;72AU:6Oc9W<2Z:-FgCaY7[E9[61_P,R
VR[E30P\\T2fC4P[FNA74<H>_39+Ye^_+c[X9_#[5:f;S/fG7#01WTeI3V2-SM5]
Mg7:E4@eaL(f(U?2AIR;?AF>D#AI4@&-DB89&\=-[[T+@e<fP]KIH/;adX13,;JC
Id9,-CON25D0.J&SOU760XGDWYK5R-UY&Z5F6G0>.1C)6H>8I^6KB;.cg?6E?5BJ
3AE,=]5@/+cAYN#D]e7[S-.WER)fW)A/NcN9R^9VTM6G7G\C8dZG71PG/2_I(+Ca
LAD9c_M[O(dOL0^R9<D17<S:4U4@#0gg1\:G=TA+3C-#J;Mee6\WC(]DfF75T4TP
27#\4I#=.faX+Q,<#MDG>9G^R?T=7gIY)@_022ea7DdP2LL#,6We>3O<J27V-NN<
3TML7F^92:O2\HT86,-DF/YDEG.a1L^(XH-e_1#V]#g[^VXJ()OV>-F6BbN]14e.
:gd08DC;;#Y9P681;[Ib5gQZ4gH.#MNXga)2@F\cFQ,&gDDN^+:NECXSY&.ZRZbH
,G\Z/ME+fc<)5AW>Nf>B5ggbgHFAIK:8NLV:FR6SA3PR3X.4]W&2cI8U<]+fT,]H
8[b.81]-aL?\7P4W1a8X<^-<W=4O[J90e7<J;eDF:&WLg[77Hg)B+C>\Y8f3NMIC
#+fIHGEY(4JLfgT0W<QJ?\B.;7e7IJO=)1Q?WI/c#:PA0EB0ED+RcDVH7H-e1CEE
6-EdO\EMC^13IR[W:R.ESBE/f9@D>5bODN.?RgG==a#VRWWb8NfJMfDfVKcNf-6f
R_G=Y2[3B8ZH8?96?T9c];Y(J3WN3fT,ec0P]9R]6C@&[O\]A[B:^R=MPZ1_Yda)
62+<aC;571X1<H9+)OQIL</J4aR;KQVA8cLV+@[eK7@7bQ<egfBLPa9,S<62CS:G
^O-Y.=4b-7KZc\=LL,)ABf?Q?=bJaEYYAS]FYX:F:M>fcG>;-W)O)4??(Q&ebL[J
IC5ca-/cc>-.YXgf?ST.fdC]>gJ?9M-U<6HBZ2I5E7L#[K9:<TbaG#0G(L,Rca-e
<ML?[dRY3<;5@EXT0WWGc7_>SRadVUVHH\@8:O>.O+b,gZTgTQ\DY(HL\_.F.TYM
&KZ4T/beX3Q,([PN#0T.4RR6_+.D9G7RU+SKf@Me#+5+TO#L+?-K[\S6DGTTLHYB
K@T[ef\ANO+?F_Y^c4PGMV__5FOQ[C1;VH2C?60KfXg=2VK2RE+VIL,4g03eH2+<
GRGT:]V9_^A1+2<IXH&JcgeL=YW@_9HdUdV_3&NRb<V2D>,TC=D/A<IaM)ggZAcd
;&TV:Y>^Z)b@)#.+64UNT5I^U,)8?FP#FHQe<MD0&bV8Fg+MU9:1QUW@SGbAW4QY
Z4DU2XB7-aOOT\_EC3]715C3-DW3[R0d0F\GN<,-&]a2I+),Ec7>B+ZXTF1-e,P3
2B4[]>f;S8+N:2#&cF-WG1Y<cf:6^]H]K63]&0,;KD9g>b#7<SA2.G.;5>I[CN:\
(U?,E1#8?YN:bIU6MGO5.;]U\IZ48CH;0.#]G15#_4#8,E1SO8@TKeVa(R7BI@HT
MD5J#GHdESU;+((d.(>G2-&bcPM^I<Zbf+AfDD[Aed:EL?cIX0.841X3P^CBcE#d
GSE<Jc/8/X+f#@):B4(F).M^Qgc4d3,?2Kd1=XA=a&VU1II(I72]FVK:F9IP1[<A
^&+[.P]ZER/3XcdF421J:/dQb-4UBWS3+-KcZO_]I?_d#+E&L2e0+[)/V6MZb8R/
10HNDW-:YHMgdQe[Z6>a4XO[d\C2S#0dL_Y0=aLPW].XY5c@ZG^H[X/g/<Aa>VZI
)1b<,)F60#D-C&bg\I3[20OT>D9HAF4J.DIV\cP=N2.RAX,^bRB@#FK7g]fR:Jb(
BD29JS.IN9#D35@AO2:^E6=2BOMd\9Ye@\7R\Q<J:([GY,a8<4JbISI3G=SRR.6F
bU^9,>95SFQF-E<gGN56E?9D]Jf.YWb^E5fMbC2U40MEBOebA&aSL;F=I?]&aZKe
#>+Tg@]L7W:N/[)JIT791&,>.e,<&;d(E-A/d@/cRc/agWPLbF4+5ACSO=4J=Z&Q
YGHZ/+CbJ6R6gI(7RP+)-O2J=fB&,]_7375&CZ/aI7XB?U230V780+>6g/?Yd\YB
B.7a7A?O#7;;<Rd]SF>d9]G7@W.DB\;&a?,[Z8ZcE:NOP<LeH8H)=ab6&&B5-UQU
??\0^dK=?OV?1007YV-S98Y=UOY\c0RVDJ_J,E0OEXYT;IU))+7-^DW)NBdYbS;K
FF]^VKQC62YKc/F-P@/WgR@TU#8VT7W0QS[L.<82DR,5UNWNeED#&(Yg6XJ3GSUd
Rc^/?,#RdLNdP(<UQ:8DH[f&_J.E]OaeXgQV/K_B=;c2YG2/aP([[Q17,-_K^:4@
3E24U>>TBD3_LcS6+^-R9H\R?BdV1LOH[G+E+>2>SPL+dD4DdB[Zd0gZ8dC61Y?;
Md](S33=;F:W_)cgUN0;4fU^J@4c23+f/\Y;4WIg27#?[Q2W9b:;gaG,4V=>T/X;
C:bSeEW=dF^V(Vc8JZT\<99022e-0(WZO6O_Y2bZK]FC#R>dbW5)WFFLQMLg0a[G
@fdLFYaX>L\b)&LB2dNe__?0b[LB-P0BQf+/H6bABc9>)QFABYQFNGX/=e<N:E9[
301\gA>G,TMNYM<#?.G;GGXEAaAJg)L,/8g#(EeR3b2?)bg<Z1TX@6?\7#Z+/9]2
837_P.M?VbdG6Ud:NeK\,Ja:NVg;_AQWP,9+#A)f?UH5Q];2[>?<8F7]),I#OW=Z
M<e@094a[UL]&@cBP>ZA=c1fWWKI->Q[\3BQ&IGA81P>8HGWcFbSK5993;=B/V]N
ga]0=GEBQRO8@,^)>.@A6TH[ZQKDIV2d?VF)2-8N0)gb0ZU(()=5G2-=L)N&>A^X
M,H=c.9&X#_KK<:#2>O(bB<WFLHGb(&U:[KaT:3a>O#];T\dTc>XWaB/4RZdQ;-N
(O?B\<1CFF>b8eT;;-HgUVL.MBLZ^:gS::X/7<f8.&-S3?31,/1cAW^e(D,=[3R7
Ne/EeS0SL\DXY+2FFV1gZ_R&aE0GWdCZ17,XVVX2:A2VBYQ>B2-P.UCMTZaPMAQP
f(_L9JYY1f+J4;Z6EDXE&0LET0fWMeKWbNGUT:M^6cFB[f^<2;7(4I<70B7&&Y6c
L5+LET](I5N[6U&P1COZ8J]V16+V?JTJ/I@NXT8R^7LXT.,H?,gb8XB7\WdWR^R6
3^dMP&MVRRdW3]71I+RCN#bR+YYYbI1V?XYO.CE,eZ9-=2S6O#E6)9E;C\,O?,85
?OL^[9e\J^f_:[5gYIE1L5f\gXABM,W.CfLW-VF?7L/Z<&[GbOSd21dNc=S[QV1a
)AY5PETX)U0P3.-YI^Ab@3Mc^QEQC[=B?O^dW;4VE9-9W\@XE_)d@f[PgM]&8AX>
:S;,#[:Y;ALTU(F4F;fg]-C=J8]/@.Ae)N8a+W[B&aZ7,-^,)0.8NN=VPD&]=A)d
Be2Ie23EP,1N#b8g55(I7fCF;()KX1<]QSg5M;adbE@UUb49F>^U@Z@+GPaY;f3E
YWb6SPWe[)6W6?b4NSEc_.^cODN8/ZFECO]d@G.^W/ST^H#ZA@M,OgB<NSTK=N=L
#>QIQ9b;WbMLWe]#X9JQB#_<5,#QQ+W@,#M?1Z,V=XC(;2B4;X?CK^#Dd+WZ/VdH
,DN2gDdJe3NRRIQV&YGW3GVe,0a3P:G9.+LM.+gS?f)SB]#Ac;\&BU[:O:)7Jc),
H)N9_VTF,L&D/e6PT1F#A@T;._E)8AI.V<c#_H?>\\])NID7POWNU8=&<La...[3
\8bCEVd;-QTUTRZ,.O-A7X,C^Pb/[_#FL@),?IBAH)LE#E1?T.+;ETFXe0U:a3U^
a5+GW5U7F;T3gO<H_RW-4=9A/\:-00K&(9RPAM,3-4T6(,K-6gdB=e:OODbd8U]\
42(Ad0#H+B>&.A>AF-0=Aa,1G-fSKB?NS6-5C>3I4A0)+(-5H/3b,_0O-R5\#HD0
/0@=\,W,N,I[e_/a>J0^V/5dO1;)>=.;Nc4//41eX+V-+g^NFY90\,)/b5M;8Z^J
L>\/.&I[eNJL)cb8Ae;@O^A&_bO)f5\O4X1<5_5C3T>&X58:V(D1^4/aIg#g5ZcE
HA[89Q<[Rb1WT3/QGA\;M[#:\\dOMR1W-@V/<<6Jf7DXDN_+2H@bbaR+ZRFb4@N3
><(G0LDJK(H>ce:[d[/H5a<D8YX+XF-29]J@f8;^fKEIQ-OZ73d0V7C@M4\?4EQ1
MF[^C]H/MEFX^A.P).L]OM2XRF9;ae.<)&PF1#)>MWABE(4V&LHPI90JLIJc?-GX
:QAM2M;L:\\Y3Y5<d&G[M6^e),;JRbQOegd8DN2&A?0Lc_A)DSLc-Z[5;.SgP@89
MNP+SW9g&=7)\UfVW\]3/M?EW0gaA,-OK,PC>eK;QELTdd8WD\8WHO68/X-?JX3c
FY_?]^AHR,,gL3I8)>+.C5P>&1308L,._JdgMO?Db([YU24XK7>a7J8U/T-E^H4B
[+;L\8)+;=WPI=_+5Y]R4b9SL>C=YFa^NT^7WL;#.g,19#ISH7@L;ZPGDF#C/[A\
B/Q#@,^^fYCGd2RbR4>ZD+@]4_T=+bA9/NB9B[69<N=69?MUf9^A3_H4:4X-9-_F
A;^5G-Z.3,9M\,U3ASVU9[dT+,1ZX7<6d[ADeBY)+F+1<<fKVN9(URe.]b)JR6J6
YEIV\DT=GDXGRPF</5YS<>9+4+)X]RO4-gbKLEP\FP8#W10bfc\>(C&#;Og[/+<9
cgF&[;X-UEQ+/@I0GZ)8Rb>8d#VZ2)Z_CJbQLd&PW.BaZ&T@;#>HL#HC8d^Lfg5I
=KgRHC1QaGagUbEE(IL>^NAND;/3[CS08ZDgM5TOUZO3>YbWX<4H8cA7Y5:I<+KP
XAX6BG<9,QTEUeIbQP#P[Zc<7bb)<#]>O37P?0@_+6&L?^H:D?B#ROHTJ=^/UZ:E
[;\BAZ.CVQD:71I92&R^WJJgeeaA?e5X:CFU6<FJd09N6UY8QV;;-6J;0]H-1-Tb
X_X@bE:UC\2?DM/QK&TO@OXPgC/,K4451dNUFaAfC_]Z=7gd,?7Q6@Y[dZ/K5Jb.
fXYf>J#[=B2e.:H.]bG<5LALBGBZWd_;#QeCY_Ae\M&#<F#g7EIG8021cE[0d.cR
K]TQH:aT3fV28PdX1R+:IT,C&#E2=^W:68QW9J=8&\G1^P,a=1[M4R;.P3/J<aL5
F_I@#77(cZS5/Q+6b5^A)RB>X^8U&K2cDXT66K+=;-ZbT_U?d^2+D&73606KDW_#
JL;0D4\b/&//2;1#=CVR&JJUc_+GR;ReWPXHIbCXF#e5##>Cc86[KCO56]cLcT85
1;K:4Uc((-_)f9T0)G3_@eUB(NBe(K]Z0P6-1JB4@.@A145@ZW<DH89dB(_0C(A.
aD,;f<WE-8E/=HW,ST[4C0VbJCSe,N[\DJUS>HY1?RdR;?S(6J@=fAbGYWRBX][;
()>,R7Q\^:N/@eD)^#c7Dg,C<JA[D&7C^1bQOIbME>e17K\,a9@3f,VcJ+@W#QVe
&8&N)XNEc8F#Q,4/eC5Fg;57EGSKJ?[4?W;0[/He6Q)@5J@B1J.^N4GOCe^&KZNQ
g_eg[b&2?aCJDKUFU#EW]dG<A&=6VSSOP:\TUOa(8@D=Y@7_9RL#T1G3KcIN^FB=
/DZI(UB(?(c4CfePa(4W&B3^M@AD3J3Y:M#.A]&E)NF.C^E7@K\,2K1g&b11V+,X
/^U[<WcTZd./MD?.E.R[P+Fc#OY,6:)-ae9RaY<Af.Bd=MW=E-[:8)MMUf<7/;UQ
>L;<#BP4PQQa)XMg#eMK:37;]+A4U.,OPSJ2ZJX=E1/)P3Y1GMNE6E)?/9J^1G4&
A\IgDf5.2P74X\30\>?<MBbGT(HX2IR;W@<-T)6YaG+L5@3I?Kd+\9GK6&b3bL<?
4FHZLPU;]32c4F)9a45d[1AMf(AM35X#W:S0Mf,39ZR(HHB.>8fCLE#cLTc>H)RP
J75D(:eMW4E0K+JXb0X,OAQF7GNLVaccYSTL&KZ4eK,KFd(.N?(]9VUYH^b&Kd2C
d09XPH1b/a_Y4[XREd4@C0[#V_eI>^@_U&J8]QefbTYH16c95\97S^GKS[S?X7KG
f60aSL]LZgK?-<ZRW1(,DQ#dXZQ=FXQ#P5aC.GCN<4CNN@3G31Z+(]G,cUOD#-aA
GgL+5D[cIX(=Mbd=-aHeBNR9&QIMBa>#ASEK2J#+RB?L8;9KF1bV@S5-=ZYC?VYP
C0@;ZCB35?07]f-#N89(2IAg[5dXf+JNYDHD\2@XQK;#]Kga>R2;.a5365=:M&3(
#ZM\cI8]/X:I?)2/0e)WOJ#,O?KKU/.5:9C+C&12;Kf:cXeWMS9/&=fZ0>TW#a\4
H\(:(G.U#fL:PO-96JX0V89J4U_]P&2C>W;Lfd@>dB_Y0,#,XMY>GIX514-)F>^I
DZ[EHa&1^-D3FF2JB#]Ib/1?K8O=<^BbKMb.+>18(2QX34FTb>EQ/,V[#8B_\C>-
d]HDJ_Ye#C^+#UaOGdPECa5D>&@UAPN#[65^ZM(&^^ZQQL7H7RB)IIg2W(=Ab@,R
9?G(;[^8Q>A[3J<O4ZNEYDAS]8(09KYU^ea<d1XP8DT77N>.2^OOA9Bd##LDH6bA
YfWL#d?-?MM]2#e.W617GR<X2N=B)1RI,)ECOXIT;;aN,QCK9f=P7Z_=+N0W^W(L
JAJ+6XUR5Y9Q<1;g_X&3_6>.CP;FB?aD/R>d,LO8[/J\bb6)7e=YL>3;Wb4LYGWZ
bBZbW3N4QA,f.+_SC)1:Ze7cKDZ@aW:X:9.\\#XBH3WGb.A&F.SJ^C#(\K=3IbM_
@H>#H.5[I\GPaa-#B-3=-W9<5HG6A[RX/KfS98VZ[)5:NC_UB+badH4cU>TaAB+4
3G02^@?TCGT1dM-/#eaMILIJ2+Z1fa@VP-)f]3/?c1PB80548Ae/?CVCQ<9,@LR\
,?:O4I++[cJ:fE,fBCFe#F/VKSJ^dFY,e@0,_KJ8(NE^\^fGUP^CUb)EZ02N.[+J
EAI,-,?4cRI^X=U1(HY6f;,(;H-\[JN)MM6c5=U7IWAJZY:BM\T61OJ@@DMWWTH1
4W8cbGUGA]aFAX4VHJQ5\T_Hfe<LE-.YJKB?]P<0)5^HGc8ALb8a>V<(D48GEVd9
2#T=S4B]26HOPA@c7NX92c,2Pe;.5/YWc0X]GG8/X;W]882V2Q_(HTH6,(8Tg5I(
Z>8.P6U+8\A:,DM_BH<G4_<a1_L;dP<;#QED;aX4gB)1PBH+2=/)W[1HSgE\N+EM
d0ReZWC\e@Y(</]8?2_WGa3#aT-V79C,Q:E#aB/C>gbT0+?]dc75[WB-I0MOdLZJ
X/dXS#)g/C=M>Sf#.6J64(fQ+ZI<<@X/.fHG(&\V7WE70.@QD:9_R4VKPb#cbf;9
^)TB7SWX5UAM6/f8)D=IPe\IVWRb2)Q\+I4cNZZBZ5Fg_5XP<DAJ?R98]AdBY<1<
KM2AQ/gS7O>:7@L5aW\+H6\SB68L(b9V_Q5d7Q_V?BC27f(e@9c>_Q\H\(8X^b^:
KIabCaK5^M[MV/@fJ>](W4gER;,S^gdK9,P#1a^ed;HOLg?ff2d4+(OU.K^\6X+P
T1,P=CKTR,c:9.ALP1\G/Bb<-/XR09NR>[[=fbL^;CVCTSZg47Y6UTbDC6OM(1YI
G15ee7/]H\PHNR/S(e(=ZE3&\(\+4PeL6YcTP>GNcT9>,+X\bFY\Y3E^?BC?K+PU
ZXa&^NN,CH.T=#P&W^c5]@^a54EPSGeU]/JOU\9D<TNRV6g1B=:D7CYC[.Y-3A65
39+Q4AI0f;K;HF.-F/#QMd7=TU_PNL.[XMHbI]S.f[<@S\WLNg6)KMHe?+M9.PS<
)gZg;6DY)[3P4cA\JeJdGbC_P_eU<Q],?P.S70F<H+L/KH[VF;/DGa=LS.)9.H6Z
g,)04G.O-2:M,NOIe^Rf-R?-g2g]c0PAG-P&:ZEaeX<<9(G_Y/Y4I[G#C-Y1H;L=
S47[>)E8H.VTJdRf_.X<>:IFKR_?7XRMGa>K@)E<Q2&>:PCJdc)XeGM,-_S=KV\?
6(3:4=[L3DBE&cYT0)G#UT2V@3PE@O0&:ZH&HXB+XfUdKU&\^,SBUb/=ebRG;](Z
^NQZZ@,=BgI-3P.g\>fM)AGb84eV6D,^5K=1f?^[Z<&GGDF\F&]CHG22S/:.dWgV
]Oe,e#.ebPQ(8B8)?fA,=?XW,f79:&^0\P:#PS,+#@UUYE96ZZ3AYN-MMFR56.XT
K1+<D-9:cBY90Z2ed7[RbUNM[4^P6W]MY.B_+^Q/_@1AP88E+N<XJH\\1#M/.[NW
>UB5=(M3XYa)3?6beD81eQ.:LF]^R-0.#K=JL^FKA_-FR36?,PQ6J4[ERW=\c(0b
:NYKc1:7eH4fc4UF(4<bZ;2;Z?[@e\1W1XeGN/R9G4S^DKH=E-a@dBLUNdfY9E&6
PLa:Pd#\^TC7&LZM,81D;+@g\:gXT:?TR5V^X9BM#F[62(MbD.,f+;CL@S.&//F2
2ATH.M.S3GYDE0HY-);Y1RVDY)1??WEV>H^(U17)05eFXW,8EI76H]+UAMJP6JdX
7):c#W;.,/bLeP^4R6d5cSeX(:[c&U)(&UKKc_b7c/ULA^BIgX?3.,RRY)ZT<ZUb
<d0B13FWXY-]6P:S#6g_eN.1R1aBb\>^Y@>dL4HO<2&)U+Fc8Tg>UA[RJA47B8.8
\&1H_<(A]25<ec5b4LUBIM7g5+NTGUJ>)O(95e-VTBK(A)1X(IXaF7aLRTCb_d1X
f#3?2#<CJJSV_Y9I?,<@+-1\:OcW(_BVI3Q+_V<IWKcg[=aY-(#5A^KJ:5:[_b@5
N>SI)-SJ]:X91L>LZ@PY6W7OM:H[ABbJB7^-YVG&3MF<WAMS<Z=8.d4ggORJ)7g2
R,VeBWO@[BT)g2LF-dYARcd84(G0=0cDJ+KO]L//]RNeOX_R:eS/RRU(9<a>JDM+
<Z-Be0H_BadJN)[O,=X-5G3)c[OZND^7I&N3gGT#(0P,P[((P4\3D)0g4LaH?gYR
4=BY8NP/^;737-,1Vf9BP-?DJ-LW@RQY2<(,F=Y)C1SBc0E&2>S7+A-)\?BYN#8^
P>VYE(ZLQ;OQ4e6TWLDe/3RP5UQ1^<FU,7UQ&)6;[<2W1GV_62@T7L-SIQ[S],6\
S2H7;J)T96@fRLLgT&2U8ad84@G:Y]AVW+EVS4TGEGc:0(g99WePU?b[aEFc?E]T
SgLUR@1TF2.A)GFOJ+C?cabB0fA_N0T)W5FEM#+7<8XXB?WFXE5V9]Ze7UH:OfDA
N\-DF@6UXX<X9bEIL4V5357BX=S_CI#=70D_0Xeb/@CT3\T[e,HS711/e9Z>X4f)
PfJdJE<ba]^Wg3B[=aW@B&<B^VdY7e+<^,?J]eaDF)LC?D>^\4H&a^:5CS&0#Z=0
T>@1P>6K:O7TJA)R5:&B:WJWeL;&&IaJ4H+12d>2+D5X0:<O99+X7O@U_8-Q)aSW
e@SBDZgAMPQ&Z]F\87cb_LMUfQ+8dV04+#T=S^c9P0O<WZE[T^5A).>TA<?W2CR1
(b:8Z@8L)Q?V-9#)J8<?5g4[0-KW.K;@^_Ye69-,X#VL_#;)KT/O-b4MY9@#H9#F
IB^A?aR?6Mb)(>)@b.=0CI(f7bEN-\^MeDUBJ+c(UIS1Mae27,AF#5G2\_/]KM:V
9gTRdY8T?S/Y.ND2N8P>QW&+X;(W<H,QLH/3eT7c4b#=bQ^c@[)&,Z#ZI&X4MG>=
Y?JW:3P^fW/7OT@e^cWLZNcRYA<b(G=[[gNAX]RU<868T):2:)U[0c3^S^[B\a#;
TU8821<?d.He;b==VP.732#6ZBUJ)O]-7S>B@SJ^\MTLd<Mg)>(EN+NJY0c#]dV6
X,RU5JU0MQfI(5&/Hf@-c>eafZV4\E_H(ea>3W/8X^0=I;?8)1QVYDF&7_L4./W?
?,P4W;C5fL[>;H-e2M>)&-.@KXIC@1]G7RXc<+Ue#X,&:=M90a5K+79+4,SX/AXQ
cZWPG/B]_2&^QV<;P00Q;O9BB[7);ZDI9,DGcB1U-/b2V)#7YQCG<:c]H9IF@6<H
WO&YJe\BG<)_FVAHZ/-2_3#0f0<eVO2QD;[K/>(WN(\KdJ(@=KTJC\J)U.7:Zc\Y
+Na5dOILF#bI]3#AffB5Y5<^1.aR9F[:3Z/03.aZffO^2d886CJ4]b(&dGO/+Ug(
D3:NB8_dQN2/a<FL70.6][OCVZ?N;^LWg0eA-]QLP05..[RNLDUZ\)<RCOL=BCK:
S]2;LY#1B7=H4VB81<3.2)Y1X,#DQ8.8Ngc=-Z^/\3d(6Zg6EO[IYAgBVHC#dS)9
BAgUc>R2bP4MU.=@d+<GO?(?#;cRUQ?.F31U05GGNRSN<GTB@+DC.FZ)@8-TS?^;
:DV3KgcTY1;02):#FHO3R6TfYGF(OT,1b(gK,d2<CPQRP[<I\0GUW3?<O7b_[?).
Q-O-?Gb__QD&F[W,[[<RXe\#EYQR1P_M\5G4Z.XS.eG-Ha_C91W4JNM^+1BR1XY#
c>@KQgY.e2S@S?;FH.KZg-MEe6,MLc\.@EfHQ&cdg?cPc)(21M\LDGg#_cCdI;=V
U)c0I7Y=[VEBLWO,-IW@13[=XXf]3f?8EgO8+462&EfCNYgTP^#27;3cJcff5?fW
aBYMd0\@dbO>gaEQ;_&3_V9=#Rc3T>fBA>Jg0c<8SU[?SJ4(K#ZbNZR//\3Y[B)/
Y#RV<0\.f_;F1-9]+73>C^YSQNJ;6U=^)54-;bST:.QVN?2CPg6\gPJRQ/@6VY>e
X01A0G-9;QK8(97H)BdD_P&,g6T:cgLY@M<_@3_5CaONG28)67.1R#TeL/d.T,g8
+a67^XaK=E.Le+?.:b-:B:8.C9(D9R5Y#0R9N9^&(VF_06+:8@L?4PDI#bg^]O)W
M8NPV9J[)U&#JO5X_:P^@&D?#LIEW./306+KU0Y7T[<BF>D>RM-)fd@V124[a^#T
;5DMQDCHe#SQ3/GZZJB\[c^1O,\:bYH)P+52?A9:7Z?E&[<,@7_Ia=\8a30K07Ud
\_/PTWVZ&<X2&N7Z#1@_]W_QK]J</2J(g.?,fCWH<TDP@eBS]TJ@F,V23YbdM1V?
Ec@b0U[fS@U.V^]db=>STYSMNgEgI47c-#6,_,G?bD7QffX(d;OK8#6@=TTS?E;M
J?80/I)0,9?3f:QbX][M0UQM9E4&E.[PX>KHL9LU\T+FI>Q5G2a10+5PKOLX7E^=
3HO8-3bI=WS.HUO1YH#YQeSI\L,AFODFK0S3>O]N5fI9@g0NHZ^+Ld+^;&K_5G;P
P7TH2-XQ;H.VZFabPDP;=-=\Ya#>9XdB0[4eQf3YHG-1NO(P;eC/SN;MXY:,VW@^
4Z\@SE+B+HC,K@cW<1MNZa_FYS18(E>T)LVaQ)eG-\aS77HFSfJKDXO.7XUFCE#A
g:&)\_\]:43Hf/P@PVAbScE.]>@(2];?DQQ>,5c3fbbXRLcd8D;eNgKVVf=HP?J-
MS;:=4A]17gOJ4HKV](ff?J:/NbC&FHB?#BHOW0aJ</SF&E490dg)N]S5:fg.IX@
7\A@_>^f0(I,8&>#UH?>K]]d6IdX&)^G+QH#=<ZXYH)(MUKP9CC\GP:[4d-5WLEL
T00&+^\EcNIK?B_YS5aaN+&N8Y0(G.GFaacJaSd4d+[N?VKE(UKHB?DAO=c)L=,Q
dP_#+aC6^>L.BD#N?9(bSN<c?>E,<-#^F@_5+M[KccY3::>_-WZf:SZGb_Ha+PT8
Qg-ZLW&6SaIdT1:WSHf;6E)g56,UG/Ef9WJ#N,>H3M@]dL)>PK,\c(#OHL93TOa9
HU:DQ?-aF62^[_I<@^C_8e9/<X;d3@/0E(YGGQT@MAQ69d+<?RD&bS0/^g7;U6NY
Z7I\=J6#cV<Fe.2fV@E4#ZD38)f=ZP=C\/9+OX]gGLUZPJV@WUL6AY5E1_Y[R6UG
X3ER81Y0;-ZC8I92IR_LTL>a<K+JgaL84Q:8\_>JMLC+6(-G\>HFSS^Q;:c8X<J0
X1P/0]RIaD^9>Hd;[e#J?KZG\;Q=Ue5>U8D]dAZ+P1?.XcE:=/3aQ\Y,8\H5)C<6
<,TDBPc.V;+KP@PBSL\O_8V=[:g&:4Oa53D@fGfTbC?MWbQ@M34?cZP7aD6?5CUf
-8RdWA_:-P:097:.P,JTDZM^WK[).BDL<;8ESA:GPa\F73&DSJV9_Z@5DJW&UZ/#
-1NIUQ^NU==3Ag7O\>^\GO98E+-@>RU3-K+PWH1?PFS+7>I.L)Lf].Qgg.ZE;X4D
.eO;&D.EEAgZ[MB\WP2PRFd/^VJGQ=c0bS/OYYPX#f35<@I>PGODQe<gWbSEZ]Ha
cd>8;>4NeREa=#g.KCNO06M=e<L?)/SNG[BT6b\<P&3ITG7&3VA_+#9(6g1#]D#=
K;:g&IB/37e)YV/:?)cI&R40SagM=O<0:@L>]-31V>/d/R@]:gbIb-9=U2]_Ta2A
POZN3AX;UZM(>&S)BC#J+2\YfbC.5Mf.UD4=5AN[a.=0]T-DRf1;,AK.6d);B;IG
I)S(^1_LE9cS@P1<^gI((0F<ONR0g\+E2S(+6U=Ng/I6D=9<eLO,S?e]DH^[\&2L
]1.68cf@>A\I7,35C7L\#-HD\AJRC?DWMAMFgeG=IfM9[+BgEK)FbH:.H4(,9XN1
#M7)gLQ8>_+ePVJMXg#8A82UUb&=#/9BM&R@CWDJCGR94;BSdUVge2J93g=b2KT?
#UE7Oa)cXZd6I(W]\LN(CMX=3AR,>g_EZ6?QVOTFeWCCB1&G&JM2G7/#X64OHR+6
/W7ED[Wc>N;[IRC@a8/S0U?.=9-5X]Q=X=AA&Yb-BGWX+_PFO0VU1eS661bV>DFM
7<H#?56g&a2TO-(/>1#=c/aP9NO9_U5V[++D;S&28b;F3(,8S:MQ&FI)?C8E/8^_
A6;D8K4OS<#dKZP#\7@EGVWIHQ(]GJ;.I2OKDNf2b82D_K=E8M77+LQRH;2RS_&P
G(A+&TcU=8BVTUQF0=.fg4[KBbdA^+WC8\D-=#8E<.ZT45#&g&ZF?NB+8e5@c0Q7
OC(1>02Q^+TR&<[AG>K3MIDD0UNQPb^VSTQ;MOSX#&e?R1C2?c2>7KMc4JQ_d9LK
98SJ#8#;&Ra_6d]SU]ZPATM,W6Z5#b0\^3\:b]C(^QZ[MVWEb/VbN0f<D^46R2-V
O,#-6J5/9G2?KbFVBeD^=aC2AD8McJG<ZNH=U[MM#^,Ud3DA=&&bV1\RMVF,7;EB
Y&aB1cga0R<-<X&-bDb[MQQP87HSLg+FD7XE2IS(2QL,?[3;<EP)E?M^]UC8DYe]
]]ac)MR(Jd@BAJB&1UB[=6+A/Q8IQY>N0VU385D[(,<&8H)A>,GcF?KHV+U/:S0W
>5-_@;3Se5@7>@[C>5D4cc8eC_>YWa4bI#8P2,I#^BMU[8>a]gJ6O<7BC3Z2QWV.
;^3SV]2Q6K3MLTZBWKH0EW2>+4HbPY1C4(Q+(RPWEO4NE>+AVG&/)5<-BX<Z9GFL
@.3-WKQDC&Ab7a5ON7Z&.Ye].;-A]C5f2EQQ-beX^fH-LF)8/,@=2=cE9J=3ZO^.
@DIUE#Sc]JUOLCf_V(YOU(8T:g(9EX?PGSFB\OUWE1<+Z;9OKG#;NMLI#HR^DRL3
C]IFUS75;4/I7)E8;Ig=?b2ZXHK\V(AaL/5cMZ.Ga4P,I<EeX2De,;?dX\)&XAFO
IQV:LdOQ?g_fQC@Z,]8[dBX8P]I)JV2<S)014gRc>N-/^@QZa2cRb/bFV4K9BWfW
^P#CUI5^[6OW6;NLPe9MU5>#Sa520G\Ecb1SR.OQVX)_,DI_+a1KYH4b,2EL_IAV
HN]?#JSB5fcK8fL2Q^([f@;W_c>L(5ETEXL)H2WJN1T=?2<#7:3\(@LIe35:4KSX
[?,1S7/gEB;d:HX[6FDJIM_N10DD&,Yg6[M@#&+)#N8C1U2A4;PQDJBaA?HDR90#
g,2#DN6<Be4>O)6/eb5W[HH/Sd20N>1[4J(4;,2A4GQcKdQ=fM#>DM>.gCgb^#[X
=I<;\,-&6UHfJLA6.B^QbTT8].LGHV<OKP@a.ZPC+_@OUJ7K1^(;,)fgZbaOTK07
)d8:A2\]4V(_a9/_+R::STRd3]8S:6&/^3fNUSf+BY-])F#BeDW8=U6YfX#?HNS/
KQU7UcL]ECU>c;eFKCYW2aZAFLNP6C4X]C+.RJM\cWObTO]DcFDfC<c^._2+I721
:.=)cVQ599)5#ZFea/eG8TDHU^Y+_Mg2><@caD2K4c1M>N(0g9-1PSIeSb]=Q+L9
DJ2X2TX-MMaY[]SKWA8MJPcf1bZ1A^F@0)H(;gg:]+6T<I1UEd[)db2]J=RJ):P@
Bb@fF/;0,V(8.f3Z5)H.<bO&=#5(;H6)c\;IMaGP6DHb7,]V[[NIb-ZL.-1F->N]
CX[VF[Q@20A4;(=T>@U/CY=0g8>X73f-^CY-[,1&ccQ0fKIJFE9C.C#6c75@)XKd
B_b64ECMCVeJS2)Y+34b=:0:)-@D<A_ce)#PPVScV)C93[c>X3a=\?YF]@G67:Y6
6b.2La.C[)]>#Me0F5CW]O[g64JS.4<f<gIff8^DUTCa=]T66?Yaf3Q7PJJ[38W@
GZZ,<FUD-FP@&J^P.P,VP0,cSfaU]R9XdTCJS9<J>Fa?b^[2,<K6R#90@>KIT?0e
I8LKSVKeHFDF4R)QEJfK+f8U;)NV70A(CCQHW)6>9a(4J8MOQT[V5[e5MZT9#0\c
EWc+1=Xb8O_3>f58_VAGf-ED,]1,Ce+:[3GAKRVaI5:QNB:FBZMaHJDY5@Q4@BS0
KMNN<#AcKEM<BP>7\IeB6TQg]9PJD0R0:+^><D\SHc5FTF(T9ATO#S2ZP@FZ/,QT
S_R\]B8eRY,6B^LEKbb?dRF,N3M0T&\cFa5F;Zc]Q0&.YU9Q4Z:-=EaKAZTUEM+.
<1YQN8aE,-F]H=MC2)K1SaC>G^JXXHJ>f.R#P,/_F+_D]\2-W\[f8H4VB^g\FKJ^
Y<2/6,Cd#LW0F,=]Y0;1JX+N(HLeW&6EZA2<HfLJ@<W&P?b(.20Ae7cX=)R^Z3Nc
<W.\4;d(2KW]?_0]QSb:;Y[FX.dbG:a].1LNIHKd5O.]6#a1dQLA#2C[QfY//CKX
X<-_\R?<\]J;[?5V0?W;:.&,Ke6bf9/caHd=)\O>)J8)W1O&)/&SU+6H;e/1O3g_
<GZ;-.W6?HgBVU:#?-:XdY<W5f/b:1-XYbL?W6a+]^@],cN?NPJ38U_UC:0MH2Y:
C2S=fL?,04F1Aa9]J>Q<XCJPOSbDRB18YJ[HE(S_(d;SA2+3_.#?M/53g^4gCT,B
/b\(e7A,L05??E/7[<f3&AJ1MCSD5[.H(CP6Z<J1C?N^QC:_8++=LAAQPfHNJ#>.
8Z#I>.B@Z#.MDN)O)OA:,=ED;f?.L25@K.7&(E@X&V7Qg]3K2H-<5WR:)A1af5\.
E0,[Ma_Q&UO]12MP7JZ5XIAPcT5Mg=1^.GF@OgLB?-[D#,e:,@-N2#7MX0[LV=\J
^8cT[].4TOIN5Wg+]SeH)Ud_K\91C9<9H><gAT;^GU8+5KPYX&?H)_YWNO[7_K5L
C\[KUH:KB>69^PHY288=WgL;@X1,L75FX;Q[4_UYK=7LQ2.S3gCOb>f&I<L)\\=;
?ERDE;K\f]cT[e<G9DY.GB]YL^>3b0WYg_E&?8?[C_cTFNDPI(,F#;aT0(1IT7(+
;7X/bJe2MYHC9B?>529/KcL?\5B6RGP&TX4K=YX/SHc)Pe@ZUOZ2WY5P(X<E28]g
\];G#aUA:8f6?a6K.WDc)?7=.N9d,LeR?GE.bFR<gVJ>M]>Z\fPeeAB15a)JA?1<
FWeX6Aa^[8/E[/9Y<<cLa4fM?cF?K:0b@-PTX63d71L29NZTB\CDc^baW2[0-G4Q
SH;:B:@gO>7GK7/BJ9ZJL8DA9&J)I(b^gaL#A9CMQQ<=CW6L(Jb1/M&,Pb6a89>0
fV\76IIb?a.8E\X86##B+c&/NKB:bAY>b<<4B<g^Ua@c1-[QP.)O=T_6\(f;CUb)
112MXB#[#FNEbE:aD4=7FS2CG(DF&g:@77FNI-1/00J3<e:bdZK7@8d^?K:<4/EH
-NJ6TTH3V,)-c[_e?P#8?65b1Y-KQ3^.-a,5d#D.gdB:O:_b?W>>EDa:V.I8ZF;P
LT6-WLN#M?;/TB:?;X6(>G.0D6]Re@0e?O7MRZ/d\(:aBC\E16+dV6==fV,51P]b
f&cF8UfZTO\1E&@aNJa.ac-_?>>70[VBFP(MHW&SYP^FKLK[46=@cX7_3TAE3S6\
<MdGEP=gCagB@AN_S&2gIaD/3.?<P4X5?YdLfW6WdEI9^W:#2=WQ3@5AGdH^20A-
4(\&?:MA_]K=fOZYO13f-7>&^e1f&2\NE[@gWec7VP][27SZXFE#<JL-(4Td0D?f
>.4_-)WTbH]f5dQ.Lc?]AO[I_5d6R@(4dEJPM<LNQ<A]+bWY+WI7CU;G0>[)\Q47
TUU6Z-\F662JFd&RPHY^L=G4VQdae#\C::&IP8D=e+:2Y__<Ae1]#]Y1NOe;S2[\
#<??;AN\\;Y6]F+dC5_#4=(#2R@Q0:Q^WN0=)2aVX_=fad^R9U=&RMBCWC&CN1LZ
Y(G3:M,]75&]6[Z&7d_BEEW2EQGLJE0\?I3EFU;QC5;]M(1X_--O:3))=YA7LXZH
020M1#Q;KCUU(FVSXNG,X3<DX-BFKBac&??SaNQQ,Pe4N/.UXN9C^P\C&Y,Qb&&@
3,0^41a&Z)AI0Mb(9_V]&XYU?\PA?NdU4+;0U.UT[7c#[Cg@,??<R0OB05:f]dT6
8=T5(A_IHOOSS4X?,N-IJ9RU2Zf3fc5^NK4US::CQ8UIOI0FCQ;_2:^2dgM;>WU7
@egU9MMD[.[EDX4SE[0JAg-GMLN)[)DO4&>=7B\[@_3(R+[5+HMQN_3N?KQ:EQ0.
=B/]7/UP2[=LM?T_Gd7+56]<_egcgW0-+[7-M1c&8]3g\7T7f,&+AJ;D>b8^Y&]1
Z,YNe\O&UZ/6DdQJ<X.)>/+b_Pd?a-S5H=e_I\86@:NLJEAJO5D3eKO5OW5b]A3V
USHW=HMC5&WRKdRM6?LK?.b;\e^RDG&Xc;MaaJ?Y#Z81^;@8XE:DM\1\/+899,>D
TY6A:^],PVRE6W.UO.Wde2YbR2G=T]_[(V5NM?d+87;R0e\(S?3#N_W>##&1JcW2
_S?[Ma].dJJQeB>f4FeS>ETROS76ABAA6R-e,<OO;,\QG\G:DM>6Og0+ZWTX5Z]I
7XC/-X,:eH,.^B;e&][?T/91U?H3DDU;9,gU-<NI4BM/#fA_0H)USI&Q771f5MV<
K[^[f/T<FQGBC:[bWcUT)Z^&fY1F(6AZK+Q#SHY@2P#O=+;[5A)5SQ:7e(e;H\YL
BF>9@&-H@;))/7UFP:Y__RJ]\#5D)H7F7aQ1(/e=[WIAIXF_-N)-ECOca/^]2L_a
9:IKM.IcXNRS^L)V1G+-JK>Ud3<?C\/J]DV8L;]643#CV&7dTMQeL^@B0,?/@8L/
g5/c?_>X+.Q2;?8Q,,)J@/LM15LX.:XFIb/f+V(:BRZf9,KW2K&X2g[,Q\@6\Lc\
>1EG22Z&MUgdL/I@]];a=CQg>ZHQW_IE(J/NUUE_;-JbHJ0]L);OWLZbDYV[J2B:
?DCd&d5D4N#F8:K+&S,a)^e[MX9-]3N4R^=bY0XfP(/R<:U(a\^B:31aR<R&P^9f
.EbTU9f@6Sa0>PbM4+5a5Q=.CWNM.5aCR(VI4T>3I+T+(N.S7afdRJ)0Rg+b@.C,
?HS/CcQZ&TRFS;B=YRG/cd1N=f+?LbT5/9Ng<1N[FQ?E_=ggZR^RQC8dWSK(=28e
RfN>bZX4M(cK0aTGY;ZfCba8UC0bcFa-()S/^fZ/K4:T:M>S-/f2&0QfW;&8_(Zd
cV6\,S&M5[_=QS@C-&A]ff\b3YA&bL2+W;:O;FY9/1bVe79Z-K2>7;W,M0CSD?CL
Gae#Ua5\.DJFZUEI3&)ZM]6RLY1NJ.<]N.ZKV8PP#)\JdH&L&1L\UEL2E=A]BK3_
>4LO3KdM\FYQ6BG?A3,BT2^>@L,PPO5X@[FcT3.ZI,eX5=VB0D89N5CA#0R5GL:9
F,-43RW4(K6./1?<,cPRV^D?@bDI8-1cQ2dAX:>OPA;AQ[-(TL5>O2<fO?V#YXEe
,g]P31L5<gUX,1+FK:-^fA<f1N;<J&PfRV_G.;+OZP5=U)&)a-M:60WU<VI&#U&4
(U0N>BR->LBT^O&)Q<<0KXCf@45&[0JRdfYS.R1[1b_5G34ZadYJVLV]Ab^1M-;)
d,8IJE_D;PA^,RJ,[7ZM0<?JQ1MbgU(7&Z4A@8<<<g<K;;,d5b1MQdd;N#b2#(@&
FHSe#V)aCQHMTVO^-_aTMXBGc._&J(_F2-69,QLC\I->6TWY&DbD17112Z9I>J05
d,9e7L7@P;Z94g7VB[J\Ie9.ANac/ICPRZS0B@\VIUS(VQYUI/L\f&SOIQ&]0Pb(
<]5\D#2>4:VDGGKT]#,gCA(FT=ga7+5Vd83S>^ZKXb<gRK<..R,(+?2]461KRc/N
A^OU.Rg\GRFDPbcEVWP7@@N.U<//VACd^O?0UMPS6YfTE+f6fXWSCBZ=+/W?\^_a
b>_V-.A=UIJaa9QR7AbWWU/>Q4SU)3a=)9I24XHdf#B_D8eb9C6b>D:.O>I6QSf7
[c/R3K)=1cbIX,6c4[<9RN-HMbG9ID[.3IVKSB4).&W(XGGN@L5/\UH]J&SAg&]2
IKC+Xc]P+L:a=RNa4J,U,JO[eGM)ERI>M>UQfS7@J+Ee)[eTYY<g].9XVQ#:LI&2
MU.0?<9C^2[2JAGb:Xa]7J4D8c.=bJ9[,3I(2IOXgbRgaZS.[a?;GSEB&:#0.XGR
[P7;#1KX35[#:S&Lb[XVBU?NKdF+646;d(/M#d?PPNY76=Oc&.9O^G7a4b:ON4Z;
?XA1,M9PHWF#?Y22+CI?9bVfg>G.bYQ/1a.a-4U][=76ZOA]AL0?#L:40H6^LTMY
I)>22H0Z6_>ON(d9#3SHJPa=&/d=+JQ6\XV8HTb#If>8A+[^_@5M/<VL#?H,GRJB
GKN0CVdYF\f;;0eBJb3?6eb+;]F>7VXb?H(_=PcZRMZ2H-.PECJXcbY5EEQJ898?
]TX34Q.;8dQXR;N_VK^(9Y52Hf[3I\E:.<Q9c0?T+_]fU0R0\[DP=R&Y5_#De\.b
b_,Q^5RKID&8@KAKg7BAe=SWJ9<]b4K-L;^4:[<aP<4]cd8,JL^FI?#R>R\g8c@D
D:VacW.IP9Y(28;/<D,,VfB<G#2+MCM,.G?>[d6[X=D6B3ES;B&7-JJQ>8#V<aXO
ac1bM?O[SHAbS1eDB9)7@-)Y/]HH(1fI/T=X@&VU2DR0Q]>4V(;J\@(@>W2a=7g8
)7MAdE[P90bJdEI+fad:1Y-<65<4gSFCB_LFa6[F-HK7(Gb5][M./XWR@GJe\DCW
G94PJJHF-2T>G-#G[a1VKf??]O-Z;&P)^,2LeaK6HXGa:+4-6Q6S?GY#YfBM0<XF
U[YdfPEc&1e5aO:]KR-/GJdCRLR9U5:Nb9RdL<0S)LcWZ=D<XUPO^UU5D2?Kb3=\
M,/LNMLPgf,IF^OO_62.0\)PGY2FR5KHAAdQ8FVAXP8]C2:H,,eXF<aW>+X9AcIW
RdT@SRV0aW4CWXBS7ZM[SX0VT[V)\P:EDR8/JFL]e&_b@S5^@XL;g^c9?TXKM_bU
7,b6b6(^3H>?,aG^OMfI0(XeIQg.H[/BK=+/_6#\Z1I=_Z\>-KL+5a\OBEbb=G7>
+W3bM]=T<1+<XQ?8f,6Q@7?JcZIZc9LeaXA);Y&4L@;7d8A^d/8A27=N+^8\,_H:
W)VWN@_J:Bg+d4Pg5;:/83T)?X+T4dN0]45>;3g)gEZRZ+LPY_0UC(LJeMddG_BV
>?]adTB^][7g;RR/,CQ8(M22g6bH/[TUbQ[5:(+6]ET@Ya]POQ/BTM]N7\LRGNIB
P1gO-JQ(dY:^)[3F]e]&5F1XfVT@0;=O[/934F[[cKf7A24WKcCD<25HIE6a7Vd2
GVY&LVc._JAf,\D7N@])[W\J0ZOZOe0LX.?+N+=G&FedZcTOOEgf8fC\\,VDTId;
c:Af.I=GE,cA04GV:d=BP#0@_;S_)Q4)UQTP_HIG3^NI,6cg]U.B)8b@/R\.<9U6
1..Cf<a,7YCb#88Pb4?)<\BXVGQ.9VaJXKA<HWECeb.4\8dSHQMHaZBaYWeaN>ag
bfS-LdFI6c7b/?g?^75M@c?&#GTaEa:QCH3+eQZW17dHL8,K>ASd8TQf7gCNALbK
MKXDS2(V2=:#PU(2BadK[,:);eOAOD43Bb=.IESO;FLP8L2@K7)J<_<3eZ+HV]Yd
43dO,45P>_WTfbU)P8=QfcNDDe#f0QD^C?6>ecbfJ>8b;?FPNVcG+JD&TIGfcb4C
]G@Y91Ld,e[[SH)]DEN8ef=LMLP5U8YUV2;A+I3,6NI(baALcZL\O2AM:/5b78]0
,a3FbOTOG12;39[E3(5[Te)Me_W?Z5#XP_R]\bXOf?fNg;7S56Wd,)(a3Q25J[Y]
F,1D]dIKcXL)(G=C8SG(5I#[>_]1^:@;C0DD],Q7YK1ZW_@?+?+]IC=eJ2:>,CO?
U+T/S91-)8NbfZ/VbAga+Z-6#QB^P+..VPfXRIdc4<X:J>&&?T7ff<QTMZ)]J)5L
QX767N#a=,O&UW)7RWg2AMc-4LP]+L=5FG-?g.SC0=e2:2&>DeQ,(g-9H;.<CM(2
f;SLgVg>bG;UR:e+UY/LK==.NO235P1FD?/1H9Q:,NO+EC?=0Q&,/DVZ.M0?CDG=
1+AAIV^-g24aZRD:<YMV.-@[Q=W]FN3=7-,B4f=.F^a2(XJ,^5B=W&U4H])HbcBZ
MQK9+2fPfOd)d[0,SN&J>T5YF21F5,aFR_MaMIR,@).eTE)M.(A8,9=Y)GdFLB#F
T>_04bIQ2c1.:=>AOW.C[a;Y@/TMJc4eC4^2d_IV)_c+]@M9/E]88]c0#2+OLBAM
SE(MB2aI3Z#4-=-K#W]2I\PC5(MI6HO8??KG8^WbaG-#)1,W8&^F[#fGT@>QW.Be
O9WSW#(-;3?[SP5SO&76L>#HXUR5\aTZI4)1TU@G13IS,9:D_V(>;ISEA3G&VcD5
d=3?[5PVHdNeD>cQE-P9WE8R(#VRT(5eeJEfegM8;;AO3/?S+)L_][d?RF+A/Q4R
NR@)[RQ\3(<5#5L==-]4<\A]GcH6UB,]U-Yg3=aGR]905C\ZKG.KMLT<.NA+K:X=
9HWW]53/a+]aPQCgFN2T(Kb/<GEC1,?SfG7P1JI(/9AR3J3c)eOH5TA3L:RT3SE[
/YObeMU)7dabETXAbDRd<A0C\LGE(D\&EZV;V>,GKN&>KN8U-g1L1LGO;9+\NU(4
YE?W[L[^H+Q<aXST<4IH9X\F:S]bYUX0#>[QZ:aa/[ZC^N[YQ9GgD2MLXXHS2(_L
<I5R8U+(:f/Z?5]b67Ee8,:/SEdB\GU\P?Z43UfWVg?b98GM6c\-fN@3dL_B./++
[5X-,:B#@[\02,V2bY,D@(TU20@HQD&@H):_\RXGV2/;OT1<H@](\:A=KRW]gN56
/<e/4fWeZe>3RTeNJ5E4>-<X+@.+3@+Z&Y&I&9V^RW/)bZN)fWea?;9)^03U\Qc8
=KR9H.cfK4Dg4/b2&XL/\RcL#@TOAYVP2,58\FY.gAf5;BQ768JR:3L1G\E76[_G
5-TJAFTT^AE=Hg@\]9R[3M?,3,&P5@\Z(GG-S,^J>[>K,@M^gE:LV\d&W/aM^B9A
d\:]#<7MVQ@[(Dg0E,eE7bL,G=PL;d>(?0]UW,d@8VRWTGfN7//_,[7JD&F_IYIb
1O?U]V2B8[NB?@eUIc9H-dS;FR;5R-ec[O2_g<NGZ4Id+Y:?^;TH_@RNb]P#J.D1
?E]K:R>.BE4<I&I3C@A5gX7[7.@RP>&\RME+#UT/FCWcG-NIE_?ZDNUHeG.X/UA>
6?90Ccf=fB+(X[2K#KC3Id.0GB[c-.;EUXMOOI9D5N+gYE&S<d:,(Xd#VSC:B4\_
WcCS8([2H>>N.9df;.V[dRC;gK#(8>YZ,;4eD/aKa;@@P(3e:09,WXAWfZS@U)<3
]daQQ7@bEc)0T^G8)X_Q7<5(,<5;&UB=(-+?A1:,32@]bZEPU7H-?:]^5TCdJ>8\
fZ9aNU6/7>R#(b@)VI1fCU16@7TfEE@01P]VD:/W86VbE;dVfUBFVMDJ+UBgM7CB
ELQ36\Q^R;O2fKac]UJ[=dW@/BKY17D.=AW2F>ELM?VXb_Qc-X]aC>P^/0T\Lf:@
g-\M5<gI;W#.2[f+?0_&W8+YLGB97=M6ZU?VN7CCJH^J:=]OMT^4S[8;H0?D?R14
M],N[^]+V39?2QC9HRJ[f)gg0XQ#D]AD,UKK3^SV^94-ag)U<#S8b)_=()DY1V-D
2-)UeX91,(M?^P:5?04\8cU89fAX_J.efU]>+7@:+DV#2f02<681b<Xd3f&H.,IJ
YAB6IVJHTP<Nag]]J,3OO7bATD?aS2X4f6;R/JIT@.C43F[RY/>K7+]8a7-daL^&
L6f2Z^62aLAA[P,;;AX8\6(g-H1U7HOfe;X-0#?B:;ADRg7<Z3+Cbae)^,8a=a>8
fG8;#)CX<g@&#)aT](U9f<4;L_K-0We6eB)==Y:JdR/7N]\XbW[\2Y?\cgfB_)A_
\GbU:]Y1R/C8GcMZ;#(OT=BV,N3ca<e8&Ka;E7VXG+J@KX/BZ0@<,Ve5NL)0T<CE
cAg@QG&)3SMZK6CgCT8MNSWRV3M/f](\A9L4fcR^M1[MFg,56/4IL^G?4P:-L6^g
/aGS@.aL/g&MJSP:=-G-,b](#Z:FZ,AVN+)UXMALcRc]Zd_(PZ/8?aY?HaV)WJbQ
2Ncg&ce+X:[55;D/GDPH@P->L=,I=9e5PJg#_<DaI7b8_<HN_a(>.\OTNCF2]=P]
<Zc3\fcCb(JC1)?I6T:=G_6OcL5@VC:\T7K7ZG=ZSK.=)/E>Ac&RE(g8CcaX#J4/
5gP\[7JVJ,A3;+(D#c,>I;:3A5@L&NZRG)LINK:Y\?H9VS/Y-)&QUe-c-(76-V(X
K#HEU7\Y=Q4Ze;L^,.JNBJ8\X69OU7G^#8Q-d)>(UPJSH-]VHfIPJGJX#Xg-[@MG
JR+WI&XSBNTN;f2;JD+5N4KG8@aOG=]61.VTICPDS_\/PYW=_Q-8KN/PgDFW3<Xc
^/#5YN-J7;V\NFO]@:P-Ab_;b?5=3Ub,b?W+]G)UQOggQe3/e42&B]O\:+153LdW
1O=REgL_<>H_@K=ZQgg0bAG;X71^\SMBWYWc]TfQP@I[RZ[<56_L\NZ((1L2=3;_
P,;H8ECQK^5_?WFE=^.[[fc#D[J&;?843T0]9OU\6:#29C_5I/+#;-??&&=Ad0V/
E0b+LXSM;WMc(-E&,K>dJ\I@:UWRGC=;YG2@UI5UTad\/HJV-)c>.b@:MM>4O7XH
6J-<MEV_a1<Pd]M\Nd^@1e\405-eV_[T[1=KE@96T1GVDa_I]WGL]N=eE-gf?4S6
CFTA4?2;@Gd]PE.UAVc,/>T][OD<UggUa\b4_C.CZX2A,B(_1MfV7BYZB2cX__N-
ZY/@NebGdLDAJP,W5.QK,KR]YS(#NFQd>4\&XQ1ICZL:@<\F9@-_3f6J4<SRK#Sf
,aCOYABVC.@QPH.G1&-3dY5/U;d/aW)2J)0#ddA@c0(LRg&1X+[SbNcR,F/LLA6a
\[BM)CV@e40)[(M<APW+(GAL^:G_Kg>^0;Ef_&3C?U]JZI4_0Rf,/_I^D\R;J5#&
DKD+5((&>ZR[TSY)HLT+IC<;[Ag[X\d0Y?_@_U/#=\N-:6EbQQ#5\T^e&[>N@#g#
fKE[&8Qf+=6O_M^.8>R:+:7S77@9<W.L^:C4#7FU=,:<6_bEM(#X3LQ^ZX)Q7XZU
@b>Eg74c4a900RNMUG8S\7UX+c-#=;/4(IYD;UeIQbMQ+P58;@W@B8QFI<SS.7RV
[\RT)VDK8T:JO\E:ab558AM5]U[fCUNFLR/(JPaK_54Z81#]21c<0W9A9GCJLTX9
24=<4EVaS>4(c[WK^\\@3D:.RQ:MR;,>ECZ4^f]fbf=:N=&?20VO?4PW0?)_c&b^
+&f?P5WT>;+3(0WVdC0AG1SSDc#?AJLJE4Q_gDX]8BK8U)]W0Y-LGc5)U9=J.>bB
5YB18A6U/)T+0K/b-EB8=E1,:g(ZG)JcNB^8^F<:PM:KZ[dK2/a7&+G)TB/\D-8]
5LS3\FCEUI3KFOR-BT;Mg+57CQJV[GfOKQ/HVH^ZXHUQ3\#U7Gd\+cP.:9)TS3L-
ITTY-=d\_U48;OF;-b]5,Jb33DX77W+]ZH>e:ceU-Ag>W>6V1A?WI0AZ#]a4.IY@
)->=(&gC@F?.gU@@3=;W/Y2eDbSYEYfeOC(/]98@&ZR,CWc]1#-cHI,eBb(8[4B4
B.-M#QQB0>63b40IK1J5S8RAH8=dVY/Y<S.3FX\d[M?B=BD)Re--GSYTPP)_+2a^
X3g0E=^QSS?3MQR7cQ>F>KP04L&P,#NK)A(M9g(-HRYb,K62,+XITPZ=RVQb(@AE
K)Q2I1V)W>ae+R10[dLf@+KFgCD=e9Cg<_<K0-:O+C=?J8ag=:GRS--]Wf._2B@d
4NNMb3eKJ/e@\M1>(DEC)U?.P54CQe8(HI3\TV^93U[,HKVVG<\&<Q:))0AWg0.@
8XU&26RTF\KD^M_/32GZG=>cV/I&RU4[R0S6-PIKW-K?)?.E:/99-f+;P)eb^#;&
_VYZQeL#ZZ<>+1</YfRK@6+C_-+Ig7dEY4gFBb_,.c5Q/NNFFRIa8b&/E,GWfa8M
.<\>-E)?PD/9A)=C]2/KYaZ.[WN-c\d([g7aKe[>D^?2TS15=#Q.cZ0EXQ6CJMQM
>cWYJ&Ie7]5[=#+d+_QMfU-[FP^Gg\)B[8BM+;6gI9,SSJQ;Fa[BJ<G07?eW#;<T
=I&Gc?B7;Q[)M4\9K75dJQ@NQ)/&GX+1,5+3eN8UbR&5@J2b^5>[=Ff#)(1/+2)V
66Ld351C0Sc[W2TSVQed+P2:VKT?@5:.JI6F]]SI&H#Oc^87I&PScNN7^c-/ZG\Z
MKMJ2[C]01W..YdYfaKC717Dg&#0+6ZOV:-b37FCW+d>D3Qb^8F)PS;aLfVZUa@&
N@&7V]a4[cT@c5_G6,<0b(d0]_T=/FHXF/(FV8Jcb/^(VJ_&8;P9HN-5WXU=#.1W
[+K&K1a?]JE)UOK,^#<BK6<,SXS3&f[YMWNNE>&g,WH-7e&?W9d7LPF8/^F?H6;[
JFQ3W2I,>,bHX=&4b?f5QBa#X=W#X>;:#(CVY[@]&LB#?a=YgD&;.0(UcRBSd:]L
>.=[C(7^/4@/E[]47]+&6C#O<^#ef:ONH91I]6>6B^D(U=agUR,W5S:M+Z,;GYR8
;1X>F_13NP(b[3bF?RA5egg6=U^Z&T@QS-GN/F@03966cgNdR4N35gW(M7VSW^[I
EO/MCJ@bH3J)Q&MFEg2#RHg1))HE,F_<HNT[E9I8X<gfA+^(#&-AG=&gHOZ/4NK.
0cLI1#T1&LLcB889_)90.IA2,A).e9DFX0YKLK.^C9Lg34-]82Re7AV_N>beT,FW
;>aQ>63K@gJRf((YW1ZMa.HA.N9]6##>BE83)AOK6L@,W/SMIVZ06W&0GKM?J:US
=a[DM0Cg,JF;C=C9W4<XN?)G2ES:\>PGFV4GSR]S0Rc1PF]_;g-_ZWW0:ZIWZD3W
9]#OC&LfZTHC,Ib8E5DGJ@H6?PF)T)Rf5c[IIc+NV2V&FeI</OJ:-2bJ@I_F(F]W
B:<<?P&FV=HP0JECK2\9MP,NC0de@>=a1e[3a(QfH1R=]1f5f,5(Ede\(e7.:T(P
9YY-/e=J?=E=6Og9a2;JWO0KGP)5(DAgVZe,8>(9=ECS=1B9e^f0#J>LY2J(058-
\LYR8)?\6K/<M,_DWO(JZOH/]I:46?3(#caP.EV5O<A-V^]]AZ/YS5gT2(IIc5Qf
&RT=]fZ^0Q417[0;dCRFYgS8:d5C[K44H^IHgBQJU?OMYHY?(T_K\E6YLPDX4bQI
dQ+e6=^1Q=AYIZTDH@Q=?<#Ac[d_+X+d7S3A]+B8#,>D71e0?L,=\/S.&Le;M0TB
-</,g,0C3[FJ>4H.#MQ&Ef;7c6#N,9U0:FIdV)85BUIL9aHfBe]#-7>N[(]@UYU1
fUSARAaabB53Bg)(AYF_IC7/XL)L1^Y,1Z,Q6bO2ZfbMT+::3.=MCM1DLVMG(27d
&I0U0-UbHSRcDe([E<;Gb:-TQD<C9C_cF_]EP19Oeb#6V[DNA/eXRNX;6TU[,3VM
QSd5F6AKf2KeB+Kf#H>5#c6S)c([2.Z]_T@E//4T<g^b@eEA)EN+Ra+HM.;GQF4;
/Y<1E7)WYdZ1A2&_Y6T\eYIQBKO?1##8ec.4PY&(+)_g>Q:?-=7&[F(G7UXV<M#I
7]\POWaD_:M4WZ?2T;Y]DHX[DNUA^=fTK6]@8(B.T4#Qaf@XW9[,e<8e90A:W82>
fR[,Jb(JU5O11=>U+1VeZgZ+c5&Y\43.70EO]O.JH@Pa&S-Lg?@eRV2YeT;b<EJ(
FGY?[Y2/?KJ3eL3.g+eZb8c&YW_7+3fFO>K@?D=M:L5\ZLF@<G6<67^6)C-8\0LE
;1ZQdcB8/[e4^^J3dL,5D>)&8eS<66WPYEG;9-:8>>]UA:19MC#eD2D)4d<_DG5V
P,S&RQT)A[@D,Q_faMZWD\(^()DK9P#WTHFQG;#9]^R-XOOb,FfCdCWE=.ASSgcK
[RZNSTOd,#WLH7eYV#;MVfAES?ZKb7Y4aR7TG@^N?R9TSbaG5P/SIJEVF<#=?R&X
Q+,>@3]TJ4<ZHH3-cL6-8#QOeOIT)(M)FWIA4&#J5S<LF\a5LU025;)FM&=K0fZC
f&6NP\A]Sa8/59/8EHOE/;:#TcM:BWKV#QH4(ggU=/V7@.(L.TDSD):;>DLeL>[7
S#PCITOI>[JTW[5(cWGEP:#@2E+X:gfKB2+)LC:70eb=GC)7c/U8LWQ4fD]@&3BM
6AgfPVd&[Y0.0/M5@?5e_cHcaKSOJ8?=:BLBf)=6c5EK-HP--;8;<#KT45?JK+4L
OCZWO8T[0?e2I&YTUg&10CJG__M.4]eB;>/W]8G2PA@f.]aFM(OQWPABC)\AfY52
J9?JH-1-X4Q#,g:Cd#CF?1W5SQ8;Oc\cCFF9C9g]Le=a_&GKR0?W/1.\8[J1DHd0
BBWCbb3109MK6+Kbd65X3aEH&R>19@OAP2:-\&aO41]59a&cX@G6IeIW3DU<0&A,
99D3.Z<;RJ2LD6a^2BY>Q;Bgc\gC,S3Q5d[>f_P=67MGd7AN)1V8KBgKGV2PHAYG
9>BWdS6gS2UQM-JVL97U[P/TAY-4/?BX7R-OaD3daJD>Q7Fd9\S?Q2I^4cF5Bb(;
/Jb/O]KU4>@5Ce:HYbP7LUIObY#+Q)1C,I,fC.-H0X[TcKVb),ZOQ>EV<[T672IB
V&gWS_aPeB-N5;-WSM5<&b@4:3:cL9VQ@EcH,J<I^YCO,Hd<_1I/L4b1L7J+Tb3:
g_4LA@45<L=(^fV,8f4UQ9(Ade0LJFB,-65Y1D.AWcT2<.[;T0)36UJ(;.21fe&I
XW=YD-Mg#-@?<KU]g0eX0BT\55;[c0Bb[f]e+#Y)C<WLVQaBa;<4;S==WQeB3LR[
8U0aRHfP,)&aG1aT[R?SUa)G]Y315@L_e)8O&\RG.G;=NcHVdEMd;;UaG>0_0&-#
SZa9bO>]b&Ig2S):Be-e4AQI-e@=Z7]O_;7LR;>ZM[K\E/=.W^^KNS>&SYd/S)+e
F^X+cI8dd)dV7]W@;&fMN^>)(5>FL:??19F34[(7IVJHI.)AU.W6Q/E9NS@.1f1S
Y87YFUP53D:-<:J_>#,0LES6@+SbE9SdS,fDN#JWH=Pg_CAb_?FVC[+a096?dQ.a
&:Yf+/5>YI?O;-d<AV[g<Y;<6K&B7-E.[0[XC5&,ZY?9NDJWc&3?4&FG.L5(1eY2
UfY\D#1)&]/_(KO/fF]RC3d(PQb;+@E&JGQa<IHQ)MWTE7N0=B.OLPU)L,ZdOE4X
2@5]M([_cVX=)S-QPY)PWf(EUW(]7,_:c3_8Wa+4Z>ZGfFMZYOb#34<5/b6BQN]K
Bd3H5FHA-MW.SM+:-O<?>])2;#NI];_:fXb1;FZfaO=/@I3AD1,P8Pe2F20<;/(;
e0b@HOac_\0LAFbC/W,RY5-R_=g-^Q+&,geU\Q8[/37N,5:Pg=+81[.[5@62RA),
#(]A1V@F:2T0CY2NE1H.N#&Z>L(F.3^^R>&B++;?P-fB4OLBe92Rca_NOVC(NPUa
Oe7[\Ib@S4eK,F)&c2a^W>--?@<-VKVEeR6SOPSe.aFQe[Y[B#Y9,/T#Ea=Y(4=9
I^VUL@]fT[E8/@/:5/_HVM-M4-&>[\/>AU+Vea?G]NO@c\UHG_dF]b8EDHa>:>9X
^]c4b97&+.RdUBB<.[ZG&bT^0ZE:Z,F;1K9^HNe44aI]B\63E:+U9PLHZ.OS.2#8
C[54gF8)?LH0U\HC#JN(EEZ[F;_N4a0E>5<4(03aObOb[[=;Zg;6K09Q9Z:65MKB
CHXY@@?&GK4-4+?O@C?OV0d-7^O_8>bLM&3:g/1BJOTgQ44H66G]-5FAEV1.Y>Kg
Z.=5M&DDM)]BR;B8g2@aBe4DeJ8XKBP+_),JU^:?F>0X->ZE,08(g8S.RF1JLI+[
M(-VAKNOJ2R\EXDC9)>2F263ce(b<B/M5O\0#2fTJ]CV](#d5<M:9:9]BX1\:]9^
Z:YKXa[RI\QZ7e<-F6ZF@f05[Y-,L71B,=<36KW)<>DNVIdE&IM\N\N8\L\VZO4T
a40bE>M0EfV/9(XZP1=PVI\O;0G51YN6/&89J>66K:0CI;X]+Y&.U3I#]3(X]?Z>
gRaWH_Rc##6f&W0<CMBO0@U>FJ9TNC<aDN8cK1R3U90Ye9L5:>IT=3YUCNG#fG,a
gH1Q3KS[UM(bbTSe0@gOFH3P[\SPeKNV&MQ^cdWN62^N/>)E4T8Z.ED7:MBD8+<\
T).=2W?MO/Z(g@T6Z5WA49[1,HXV37g5[A)W]8FIGPAZ;.94A^4X@1^0UM8^4^[3
W917A#-#HagVIU?(+D?1Q5H1\WFNX6d^<LY)S=#<<Lf&;A]fAE#D-BQaOZP1WMM]
Pd2)7NEAZdeMJ/IC#P:G]=IO:FG1C<\IL<.<b5A]+RQ9NC:Pd+YL,G;O8R+a#R&=
g_d#OI8dXQ[6g\;ZcSd?[W/O3W)eYeGB9&4f34F2F/GY;S?R4=GZN=A74G)+K<>J
b+:VWeJ+QEF^#((S^L&6]/-dL2bP8;X4W>>C\1Xc4R_542V<&Y9;VER<PQf#Xf4>
/fT3c)1D]L<F_/8a;Ye\T#6F\?P^&,(KW;RO((,_HBZ_[68NbY.UG[..@cR]_B6O
#M4O],/=PU09[TUM(X7:7314W=L3Kd?7fa5a2M_WN2LN&:/)GC-:E4]2ae_\2VO1
XW_3#DXB(&>4>+K;]TNe18;Fd:=d\F)V)c]G:BN6Z.(@Bf?]8SI-T+N,g&[)FeAF
U=[G3)/6PW57GKQ0e&_6HO6@N,GFaN-3G<6N/Z3BUeC?bOafHN)-VNUc=<3GI[(4
5TF\7>#DB/.gU[04X0DdISbZ_XK?8\^MT-H3>(R8_<T:,M/U^I.?=&4:ZY09^-+(
XGH30@;H;CYfe-M6-U+7f<(6g.K@dbMad?)A+AA1MQa1[C_)53gS;f5F)cdFg]Hd
MHEVS,UC]@+ccXc080G?5d_4U30F]-(1KMG+;g8f)&0XW.MNY;S<GV<F,:Z(fd:@
HVX<IEbIJ8#:_.KT07GGdaNET1\S>N9f70I#()VQ0QcCaecNSK5\:O_P[b:gOKCY
78W8a,M][WaH6VV&(8?[Ag5I6ET2N^6beQI]\ab:L9>_<[-OBARCZGHPeT=D.9A?
dG>>,G_fX:FfKO#X0HdFFXOWc@_7Y/B[IV0E6L]AON(\EYdS:LgY5gMB<P\-4cdB
M[+SJfa0EVN3@AN\(6E>X,a7-R@a=>cA\CM@d?dAgMX-STd9b7>??2M/Q1Z[db2b
Ya@Z(PO;9.L70,PQ^b<O@6E;[=TgYD\8&HdAa,#ER]RZ-/fcEHOJ=G>XIL&Q[\M7
HNRPH;E.KVC13UYEf8,HZZ,b=]?L+>SPcf31OGW];I6.Q@EXSLDZQLQ@e]8?B-8Y
c2FO5:_?WB)eaE[#C)1R2)+U^ZZ@.OeJ-]^-^R1TaPW>G+,BUJT\:1Be]+OAEX18
I:7.RVKba?4DSJbH7NH(\)96UZTA[Z#,b;/E)MD6-;R2V2LeISB-_;[(2bAfM#3P
G]H2PV&[DH2-:N)L\VfaVd@@7&deE[,U;17C=<1LH@7\CDT=7dc6E+T0][-8U0)H
\:B<9d/5bW1FHBdbOd2.^697KEAeg<FNJAFaNZ3\BOLL72GDa)NEb-W2eFH:daaO
,Z,.dS=)Le=5:QPeQ154g3/5V^6&WG<WQ7,UZASPN&cB/[ML#I@ZBR.g)PC.<+(=
c(#9TJMM&]:#C&(2P+_5gfHGD11OHG;B8g+bQ:0D/B6L03+e#MY+b)7ad\W1.26A
]Xb-BAA2\4X?,1LV23#^.GBg;g]=2SR][R+-F91?R;4Z8SP+cNb3<V+gcU\A]4._
a2Ob;70:-W>;3e4-\<d/FZKP5]>11eNVCF(B;O())/LO0Y08B@Oa1:=E=SX0?NGU
A1>f?^OC+(LF<\OS0[I0G:)86Y57,6G65<2QZ+?6(]Y;1(S]QVCYB4;P_RUD.G0g
6Y8Te.TP=0@YFDKX;ME1.e5fO21B>=W1GF(<[0d[0MaN\Zb.L>U([R7_KLW-dca1
<<f\Z.4GT>?,,HgD+2FKP7MX.VM):\FG7X(,W+9We_D]I88H5O8D0Nc)2##GG<Kc
/&;f(.:0:d-VCE<OLAH/9LAUOG+8RN3g=WX0Pf<?]2?=2J?U():LEZ(RL:^c>=.+
bWM-C\,.d/T#N7:V;2>]V>FKGD0)\DGPVM7DXM/HdLR7PdKOec-@QY>?:c)0Yd,.
gAR@E@S6PM^;&I9C6a8\<Fe_=K\AcRIMF8BBB1HO0/a7Q\>()T^.6_(L68LM?A?J
d3MfJ,Id>U/c32RTE0SbG8MP=dX:))Z-3Z><4@d2_0@7<X@dKYG:_(G6Z.HWX9J0
)XTDLHcE.6^E[Z67S\&4;;Q(XdX+513g08KG4C]UGg4eaSWPNZ[+=:MQI9Pb\AFf
N^Oe9H[J[,A?-78^6^VQQ5<]&>db[/F@67?f>c;bdKPIW>3\Q(1;eWgI\];@HXGN
D[\J8PYcOD8KTVTV?#UO>4cMZ+K;T,(SK3c:V-<)<XG36DG8P][Q08e/aH_DJ#:3
_f=&P7?V\4D<=YVQV1SM]L)dRV^1[R1_6/31@,\c.Q2-c@Zb;]P+3\=d5/f-GgW+
Q?VY#^#2M#UXLc(,143bIcAKQY@=Y(V8.Q)&W&9XF0Og(Z:2@g6>)dAIZ<;XfO30
L]B6.<R,#QJ<EYg[+3=Z9F)bS9=&(HQOX]=e2O[6e1cO8:Q.Ca[+(:8E97BIHA(1
G3NbBZHa+L6c4\+Y\4>]^B]bTH>YH0<ESgWL8BXJK2EOBBQO671e6.9CB-5=:CXQ
6G5JVLDg0/U>MY3eV[YTE]#.2;cgD/^f#X?/6Z2@Z,88H_=R,bfD(?,bC:6U71>2
=S#,&E_S:L-E:;4/-J,H=/[MUCZSBIK.F5DdST;f\SMTZQC.+b/RW]55H]f)bdKO
NRK,4=dLb,9GAbN_[5UXR]FIW3N[:/B9Nd?1Z<6[a3;X/(OQZ--a,5[e7Ae:>Y(:
4H7Z,21NbZPT5@A2\J[3c4:1OQ>KdII;AZQaP4YVPRedfJ^c9U460J6Mf.-++L]8
CPOP@95A,CRH52HS-IE<(-1bMK7+O<,8_N9AW>TJRdIZYOV8C7AQ:IBJa.R0T(<J
9I0(D)3^Da=K73eB2[,B(SI_E9SAfEGS@&KeACGXGF?.Y3eJ&d1:A=@(UZU/QPSX
?M0/UA/_WD8)6aC2J3:\-UP(EdKDBd5TL&-HDB^_We>6Fe?<FMR>OLJC92<3aafb
e]VV<^fLN8\1TLH>T[fPJ_0XXBK/M1:E2_[(&NLVX(?V=?4_I(GK3_^5/>8^OcAW
931JO^@2]708UaG\_&aEZQT>.6d4\MgTQfg28GY>VJYPeVBGKf)<-.D)fUBYHZ=F
<=Ie=KFZ;J>,&5)@:MA?(f6EWSYWO-Y]LaQ>I_g>;f+:[90L@W?baZPa;/;9/T3Q
#g_P@;aB][DS94\A8C5-GUCGca?3^^2R:.NMW&Z,U(^gKA::M@0MK2W]1)]aJZb5
?Z#bKGTC+3=O3U#ab5S1=?8[VeMfLaHC=?B6OfcVYI>_[aa@QXGH()0JQ<^N@UU;
Lc9FgE/c_EU3VNQQg/W\7.(3[2c2fa\6?#MZ_ITB;gI)81K-IK()W,HSb##EXDL<
SU8IcPSd.OIVEOK>1C3CR/a,B\L^c_KFB@gCG)L+1&R7D1DDT8g+bTU=WH4fPOR]
6^P7&/(OXZP/ab,eB_I(gS_+]=SG2=.7[9&K#LNcYE9A7M6e-P#OBHN@\=U#I&RE
aTG_F?V9I?e;d)=<JO[(-_]\Sa]ba]?0MBEMegH]\cX@ZW+JgXc7Dg#S.?>BO#\G
6d(HHR5,>#IH#[A.F6Z)aRO]YU_D0DA,U=.@CH35^c#DGS97U1G1(-7],G^FObbF
W]B)G9IQUNI=;cS0dYI29/5S&d1aLXV:N?]VV>TZ6+Z2aCI(]F+)eP&;]#O^Fe]&
]HP[X[@&J,7WUM[6X>O;;Z[FDc;>fIKAbG&7E_f[^V2J6@caR&JQFgY5Sc^8\4H#
(:\F-RO3PPDbKaId0IaYBYC:[Yf64V/S3W=/#La&7+CJVX=<E?KP5J#+VJ\CNHH-
GWL4)_ac2^[c]adYYgB]DCTEY45S)(J87VYMefDD+>.IQ21UUNL7P)IQ</X14>Kg
4&8gPK)CE15L\gF#?U=9a:L)2(6SROUR3-,,=KbU#@&D>/J)<e22Hd3?L+,H#QV/
03&QaJE23LA8-<DZbG>6P;_deT7@N,X#RSWR\TIWF6L_Wb(313@-5(7.FK0>:-#E
e:W(1b]@KO\Qc0LSR#;8<MF4<=Y3#1bRXO2]0PKS,2CYL3<X+[3-FVHL5g\H+3\<
T(D=AK,I^<\dGQ<^:9/[7:7/Oa:45H\ZQ/:+8/20C.:/JO@A_a7@59e?O0R-<X+J
f[NOUW[LJeM,&H./?&\(6[6(bSA,g^_M<G+E^C?g\6MTP.WcWH9E-c32#AU,EN=?
XV4)7<B)C?H_KNY\LRC.PeEY&afD\O(ITS7M94S9TFHaIKKE67+@(D-GG4KN)C1K
P5FELIHY844SLNN3(fbOY2VKB7>O_@C?:OKY)O[26QN(:(Y&3)[S5>^;R)_UdRA+
6GJFVO=A;//58VA0(12/V0ES+e?>LY6V>94e<SPZc-F1^cdC#aff1fWW-=<65eAd
Q5761?eV./52cA;eN0X8#>X00-5.,Q>:SVZ7cNbG8G##7\LI?Xf9N8N;K,\eKR/0
AA[LBfBIN=RT8bDV=Ja94Y<&KZ>LINNf1FS]B=\AG>=X2_8M0^E57\R:TK9X)^cJ
dQNE)U^W9(8OS/R(+ILRN<+DBdJXXQbJY/E3,9=N1M0/=\0V7Tb/)[6U<bgcd=Qg
2fabC-JTP7>]_Sd54/QP30Wd.a]\YP2V6DWWV9,9R:[(I+6U@E5\?-4S[]Jed[@d
Z+La:2C6CVCM17:FV11R=._S9fRfeeX)#,U(d+=E^FM)@gKQZ<S;-22M46ZW&D>&
-#[XU?=T)5T.[aS67_aM3bM.Uf+efDU55#;6;07dIL15@5HUgdfK?c7aG-cRV8H5
=3bb69UMcZ&DGcc4B\_6I3>4RRN@&CX8P)c]:U0W^RL4cGU96EM--:_RXI5Ee,b8
N(1,W0\Z0YAg6IJ56J=JH&I]\M#=0H:C#1Q([+U&8VQ?D+E\\,a9b]CR)PCb<HGg
N17[\7(N,)Jc)IULAPBK:>8?c8G]c.\VQ1-Y\:6d1FCfFcBaKE>VB5PBcE@K36TZ
cYE5<2V&2\]FS&f3ff-g(3ZO/[GgW27#ZTY#1b_ATB<4GbC(EccRQ0&\ag_F=F,0
b1B7RV4bf=,fZ7TDT;SLb/SX>)]\FAQ>W5NC8Q,Z2X+a6B>YYIe1G-5XK4L&Y_8d
Pc5AA@\@36V10S6,dXBX(W+VD6=32C(Mfc/e75U^D<N=EK)]VV[CRKQXO-N#M<Ob
@T3D-G@PX6eI-^cY_E/W82S+beA,W:H8OGb_@6T(OCKfS_Q/N#Zc6;RE_(9BL^YW
/VOg[-O[^g.eDQXgE[@FEN8^;6\JM;(CC7>2+P+-#O1;?@Kg9<J[7d^V+Q)6[J^K
#QALE3PfSfK:RSZNKCW4#W=)KB0e;[F;2O=(NFdf0fRBYX806?Hb54.aE[L0d8Qc
R^I>IALP#NW;9NO2]0N?AEa5)LN&@0ea]O/\dDVdOb6=./P?.1N7M-R+.;B5F<G[
9SWB>L8>9S2W=<BIOF<^-2Q=>;0+R1:J),a0X32XB:g)B\PD.S/;gJ&,CeI\g(08
Od_V;[.PB=\3>T9/YZT6ScNX>7EBc9X+DM-K<YMaAIMX.8cGVQ345Q1Q30N5ab./
Le&WJ^<I0G/:ISNaR4#4+NcOL&cI_TF_BLOC5/+_B,IbfRfM2K]E2WO<_CL\IRT7
Of5N\>ZF-DQ?VEZNW)FcU#V7C1L#O/6DQ?S^>+(bd#\>NVB8f81)a]D9_1LWVfNa
T:;R@g66#@.;2D:90\@D#XbO?L+I;4H^62I9#V9WdP>;=AXBO^GRDVMXe^REDFSI
N3O((86^4+_F63<9/;;,QXDPgeD6@5Q:b^Q^Ua6?.J#35PU,K@D^ZL8D),XS+XTL
=_\:-A4>GA3C?XC96KI9(G/dbJ8>62(2,=92UaJ&0I+e3?Q)?I(83G8A6[SV(T\T
GPcFMZGMd[VB@_BC18_^73BH^MJ07+K8__PK_AaaTEgb;8NVRWW?>b10;T13MZgF
Y5#8)+]?[EG^3AHgIM3f2QD2^;ZDVYYB74[<-C/b&dML=?=;@@8MX[L^RWT4<.AF
RJS84SD)1<F^4N#X29C6D8][?3[HfUf_1LI9N&b31AUFL7)_c.AQaVF_O3^R6QQ&
FO79UN&MF&([\(1@SZI</[VD=WOT9gI?aJ?5fAbG>f?;#MQL@BLK4a3U<W0XE9R;
#[=@+f/Gb1\1XM+fW1/X0=N\C+fE1OcZZQIS<fb[[N>a6a:EPC3C;]0cPPO;NK_8
4;^B]f4#4<O1d-PB-YBS5(Y^13N>J0gY<f\;31/R[Z/1U_X_7W4Y><C-KcMX5d:-
^IXKgGP:-W]C/5c9aE;+\R.+[NKA_)c=C.(b8OS&B\?_Q-,OQaSJ0(CC;D;X0(JI
(JVS=_60I_VI]5e93U[b[./Z([H((-><:)4DeWRNTdKW92eN#GN2Pf1NYR+F?_c]
fPLC1)D82#(E_R(9Z41@Db1^/<Sa6_=;P/IK-PT#P=gaW85PdT,gN/]:IJZ?/H>U
-Hb,I6Q6HR:)cIR#O>CFFCYHJ239K<#GT#A_4fKf\EI2Z.UR?[24^+VW39+U#]U2
FKd^>F.QAHC7=U^fZ<29X[W^@IULIdW<Q\LL6K8@:Fg\c>^>=:R@]dd<3Ic>B4:C
?@W@GTHOAF345\0WHfEd/JeI<J?FW/JTcL?RTZ:<VD:BAdG3;86T,YI]50-?E9Z\
Af7@dOJ9,N5?0b38HVB>7+>B1=ffY>T7X3P.@+(U[E,@][.CA])L<d4F3^C^1H41
c33<XW:[Z+6C/PSb[VT-E^(_e-Y-W#@eDUH=/.a#_5G=f2GCX)Y/&\OXH]T^6>QN
QYa4Jb6MK94^PQO#I,AN)^f85VAV#]?ZD/OLQP4]=6^27]U:&=10[Xg_]<5+UDP)
P+>b[X[)6acW;J.V,8T.9OKd3/.:ZSL>2O^?Q+-[8IWaZT<^CX4g#[]E<#H1[7,f
>AJO[6\VUKafR;Y-)N#.+;B\>B>5@UF1>V93)M,JCBE41R#=RI)g3A#O+8a:F??5
7G&5F.(P\Q#=b)27G9fg(;V]7+8DE,CPSY]MSSge0d8I)SG(#NeQ0U@Sgf4/5DL-
(L\GNgG/&JEH(.e7LM7^PPT2=TPg#8aEe_f/JOQJX?)77A7B7C18K0UD1(C_a<05
3=U(^S]WH;3?fR.PP1TVc#72@-acB;;fXRCJfA]O[F:I-1TQYd##LQ^&b15,9R)>
9ObJ6)ADN&=C=;Oa+]gNfIN)1XFeK-_.SQ)K&aEV,<983Y:IRJ&dN(;9feGE3#WC
D6NVETaEd]^TO=P.OdDC\<;fc,B+RdZ52P<gg7+G(=VS6\MeJe+KDHg+\)QdQJd\
(LGIa1DZ(18d29VV4YYHO:D]9&_/2GY#DNe,#T9&(L9,Y,]0AcALO_^I;M]5.L=2
G\O=g35d#Ee<4YaBc#&:c.@Lea_ZG,I5MM7&5#ULB7L>=BQf\6HVDK<P\^g^,339
bQdL@OSX(#/f3,g]6=e4:\?F5,0/MPMBPP_-^<g(.S;3#8269M9DcGRKD/0OM4][
a6-(Xd1Ta#Z<JFF[KKE+)0(/^D8ES1<4W]PCMK<V/Y=CQG5FM[/;J[NIBXYA?::I
^-+c58eWNQM=a),E.+/7eZJcTbW//FdQAA6LML6Y)G,.WR[P0L:H.H3d\5/T5OSE
SGIV-F@7&O^@H1A=a8>AI8K3Afe,.Y3Hf.>dDe#cBeKL_gdOf.#EE(HX8MbB&J[(
H/bMB[:2V_/X&4HG<C3eGBAI7V9&Y/1Vc7:]dSDAQ1C\^6:[H@F6-,3&^Jf#&IMN
\aNe[YH,9N8.IH7K=Bd:RL#AgQAg#A,,2XVDe@Qf1g2EJW&ddc<8FL3G;J)<5LC(
F+TR:D[W:]aW\G3Jc,#KL-=bL;G)\1>U.O06IVN]W&[UWT=/8bWH;AYXV#0,cd?5
6Ke^JHP[.QL3:5W^8VBH380B2V)?Q7Yb>C1.G6)4dPF7.EU^6J/ea,NA5BKI-87:
0:RL8d.NbB-4,aYAa>@(@G>^7(.))/AW1KK=6^3fZ/I>\Z.GI)Z_@@W7\2-W^MN7
/@-?@B:EZN:Z^g48g.<&4/N]2]78MReGHV_3:Z/8G[)4W;5a>eT(6F.ZPH(be-f=
]>^SK0AT<bDKDHMPdJ/]Sb(RZPJS<NDB1KTD-(=BdM&UHKCIT#)-S@HN6Y:S4bA)
cUde@Tf&6@BDZ+K1B59I>R)/TR<eU>Pe#ED3:a>0Gf5/,gN;C/\1B=<f@]FG(VDI
&/LV^M9FGI-fL.ZeA1Jd,:,@UL+=<;N2=.)^)7^CZYdCV@NfH#VQ^E26.80?([E,
M_c[ZS85-SZB.DGQfa]@,O8]1+B,_ZOH/R=&EWDYGfNX_-f-Z&R[]d?V7QCP;F;)
:5>X85aNKa_9-fF,8^\3XK#(?EP6K3a)>6E4+B2-QXD6(Q]YIN#Bc\UU]gYQ5&KF
&QKEf=\@?O[L5^_R92;HANVII5.^a]7-[IH#;CHUL@gOSC:X0\]M6bKB/\9baX)]
WD7Q280].[fFN?8CD9=-\cUE9<;Gf4P)ad1Fb&HRT/#RbAHOf3_PPEYZD4]aL#..
]W,\,V;Kb)9;R],aTPgR)60IA199.R7IaJP;C41TC=9DY;Vce#:BQaZeKXagON8#
TD#OM8\W8V(U2(=FJVS\#G^1XV1K:&;F-Z<JWWa)cN3@5b<BJ-E1#fb>A6/\44G6
[,&\M^2b]IaQ?4R)J:T97@X7a,]fLB:MVHU)C4\V0,;,28DUJ>@3O(XbE(R3M.>C
MOOeW+G3M]>ACbOaN7&0,#9=_@;++=[>N(MDe)E3V[1^TKPe;^,]0)?WaQe^DSS^
dC4MIb3>2O>cfWEX/B,TTM>f(a_@@/V6YTRfg/,GON)(bb_GP9#\;&;K5/-,8aPM
B\I7EgNVE]KA\N9[;e3.32bRTaAQ^]I#>30H)_a5V[T_9Pe+G0L21-f+,KcDT=c7
MU9g\.@d9ffM#9cW+R,USd9a=:2HV;TJT?>JcIVSUFJ,W4F[7G\K^^.\4IeE<T_&
[bMK7B;BRR1F,cOQ&ZI<6NDY9W[#_2T.T#8LZ^K2G.7]?)NREI?_186F@#&>7;eT
.)4:?A(FG9F.10Z5D^\CE>W-f>YXcY(/0U;_.OL;A8cDTWNX(V\<K:/6)X#YHT]U
a_WQLGMT=[@;DGgKJAWL9QY)=8Z9Ugc6)SA8gcPdCLH)@=)/HOVc>Q6H#\fAIUFT
H7ST9G9Y)O=dPTDK<#I;DQQN_AEf<L^B^.5W=J^H,^a@OV=\YH+U0H)C,03E152]
A+++(3G^e4.NJ(CNZO:9^IcbDI9VBb/ZgI_685\UPS^HEQbC4=dPCT)cNdNB,R0<
G>LFQM(V>W@]Sgc:<&c)SFG#S?FfK\Y7d[,S5QHY7P/6=T<<\[C.12/F4BX5\-13
E,2HfPcZ5WgDQcY#GXO^BMQ#E)YIG,ca3[=&?@N0WEZ_&FEfWVaN=19<=]3P:[e8
Fc;](.e26#<J3c#C4UL8D1(OWaKT<R5ZGM9,GXd),_T>7c:\12R^7&U5T#XbXG.^
Y4ARMbZ(;?RH,0J(=/@#85T,4N07a#<QXL]f8Ad)d6WY.2O5Fb+ZH4O54+>:4N.c
d@ID87_)?7cDD6fJQ@MEJ(IZ7d=_Y>AI+CT<EdE/K5AZQ(-BE)T#4VN\M^[c5LU1
PHa3@6P[9/eDH]W/-g<-=P:?S3U04Sc>TE_RQPS0BL^+3RaIedDeV3FVY2JK5LZ:
1f0_Y&-QB\A7H_[AK3(.Hg/:DgZ]5N(26L0Tgg#>UUC4bT+Y>e7G:bCHG#]K/M6R
Eceb188<fg:B[,5FV26PJ;J<KU]^W#1EK:9K+bSU9G/Q_8&T)YYF&QJAETcK?69?
f9W-cB7(/YS:T=2)Bg&a\f@gNJbbCDR.Na61\/(cgIW^D^J77H&2SBMb)a>:f2+@
[6=](X(O8][^]?.&L4+ED/Kca8TF1Q<4)SUNHeAEK2DQBN#J[8USK>SF?B.UX(U4
+SO9R@-8FB^L3K//50gHV^f0P5P63?J>>(^<81R#OX>6M?[3B?:MA>I=b-Gf=H6^
DNa;=/GgS+QL+ZO-(dC3-)ZV)IT)LX2#F/JeMU?7a4Pa^80CRWBRf]TN#>EP)F6^
U7T,:I[VN/HL,-<54A&ZM><@9CG06d9#&&0QYQH:E-8:08fL09?<PAMUeUC5<;X=
:ZN^J?OXa&.KQB)ER\H_4>QV7#;LV[&>[&GB(03Se_\CaBTWIFRRT6RAG>N<_RLC
9)^L2Rc]CB-1-CE-LLb>(G&aRZ:&gWUAQM<GbSLB3=Ta7WP(ZLJQEa:a;NG+V90)
]Mae34Q.eL8HdOBKTbP^SccM&(^OKed?^bH8P;V6MVLOH[6ZY,M<:+UFCEYMbU8^
-)E^68aT9gA7I]YS,S?JC7F_Aa?ZG_(YDWJV#e4KF3M+aJ-^SQdD#()fD[?(STQ&
AE@f05YE9W++GEFQRDR3YU2a,;;?/J:8L66A.=7I4f>B@][IT3\JVF77@6\aS.5?
(M-T93d[D(#g@e&0/J-:YWHB4[A/[L/F_O=D:CV\^.eg^I1W>5:;KO#bJ]2GR:K9
>b[4H,<LNb.f&ARd1/;]C2-(TLgN:f^+C-_X+U7I?HaY1#UOV@5>BF@\C;JZ5a\d
&Fc+77?&;1MdS-2SDZbS@aL-ZMM8?@@@/6;998PP[&N=5_=3f3_F\0eHC?<;bJ2C
NT(#(-JfK8?SR\N1:PZ#[RYSS/5]3]KT379HI27aSGBQ70@?RLTT70#D1+;:ZQ)=
6b+\Rb3B6>TM,5J)PXC373[RIY_E&JVeUS>P&CV;Ta6cY_[K<_^RD@E,,_CK,/SB
;6eK8=e\Se3P/gOTe9U:g5M_1UOTV.@gR6dS\0,FJI=H5)cT9OcCT-;F?4>8F/(e
X:7+0ED4bMTM&e8T/R\AXa[:X<YDB+SEE._<e/Zb;5QX1g3a]55gX;HSBOE&TS)W
dE<W<?e;_KZB[QWbd@8W=NIH@9^]2IG;JdQf]2KT>-6:-HWgG/J#Y8(]6BJDHE=Y
=/KMc]USHRX0NILX4QCQd-?U>,D/;1O68]:+?)f<:F-Z>(&]\#c@,).b^(MH/OKO
H=Q?)F2CR7YDfASH&XKCK;?;ZB:e1UaH8ZJb70?@1YYHHVM;Og<?9=]3Xb4eN;>X
-fB(b8\MI-KYB:<S]=R1G[SQV+:]9RfFXR9MN3/f-\J^;Y?cY<EJ_Ud+E)SBK.dd
c+;Z.g]=>J#,3b#):^a\;PfeFCRZ?^/(HN#eMX^S2:Q>,]_64MVTd147;Zd1?_F5
fE,YSI<QDA94(gE7=K.2Y0YTCe\I8e)?,)b],a\2[/0WA_28VO3QBc8XVX+f=?XZ
LfP&KL@<\T5ff/XB_geY7Z#7QcMeb,QY@\P\;I5ZR>[3D^;HZf;1S=RRP9e-S\M\
R./N8a)DR=F]5Q;NJ6dUJC3;\&=<?8a=HBefR7cPcgP;9Nc803R?fS+9&Ng=ff1b
f6Q9Y-?f[MGEcFQ+#39^/GS+ceM-g?W:LS0b[@+LHL8E-BE0eg.PHLAJH8+-I3G3
U8D03?@STJBC5;XNWI[aO,af+,[YCVSE6>-GW7gOAICE7d:.8&LUH0C;+3YaG0AG
7g9@g1W0B:1#8][e\S]VTEA0NaG2=Q>4(OF1JRQQZ>;Z47_TKbZ06Yae(EBCeC;6
T#f.=SQ.[94T^7QP[RSO>9QCLS+cP=#41,?IEM\#A1+OX[78.S;02<\Y]cgf>C>=
=];[K&XUT54B&(\1.CgR-ZWO?4,:73?^=3dTU_cJ?[UKCNeOC)?H)@fYX8I\<=^_
T2D_M)a<>?bRXIGd4&/HfRY9^;TfIZ(AOR;O/LXE-WUCV,N;A7acW_f07?&]7PaK
g[E?L[2.7;bNPK[ZH0I=^Me_MKR1NKNVg;b68E6W?1Z]3\:U/cJN4F80,AENdMB[
PO4N=T=701TSVE=POc\cT_NRWK9,,A&GR_+5_:USD1#PMVE6ZU,?ZC\+fWP_]QTY
BY8/B@]>(BT0JNC7-ZNN\S-K3<+JZ&P_G:GV+GWcY6=DL7&;)QgK+AEVY[79)BHV
>DP:+1@GL1W>O?H?]_D[H;gd4]:-Ge^RRQ1GMOdRX?.#/Y[QI/:7\g(<)?\45NRH
]c^^H7H3g)Z4.)4OFOV3J^@&:;+]DGJ;fU&BIE]Q@[(NZ.)G^,5_66/E?Fg?8I]I
D?RD;,+81R5egVb_H0KKU^N0N:,X-N8e-Q7(I68C+-+#,7U#HN4O6I5_]<4):DgS
AWa.SKAA2\,T_b9I=R)O2gIMMEGAHN/BaTA6LS,/Y8J+JcA<-Yc;JD?\K;NXaYb9
N,b(NfQZ7_3dCB?a6HBcBDJ2RX1P0bC/N;>0-/ZZ\Lc5EJ6dC^QTd(5INQEMBMQ2
UcM)a912/_GVK;T.B3-RV&62]6=_+)4@aZSG\;IWDA(G^I\O>fL/66aO.AV4-P:_
b=C&P-@39@Yg+X/[faMF<CfT.M^[49Ka<.IBdG=LRdYK3PMd&OYb&(D7=41-Y-#[
C)-RJ?==#Fd37CQFP7.K^TgaU2JZSbeE=:EA+:_6Nb-@WQUNL:ZUgV#Eg2#R>DgF
BU@]Og>OKB@LcFKIAJf?Q^NF>?CE)?P7H\R\#8f5Ua4>E-2\7-WJ)e)?gL5daF=-
XGNP9INQ:Y<)+IS56:QcAG02?J2:#NQ&]3DfK:;9b4#J_TZ+]G;/>gO&GBG,Q@cU
dI/UcCVfK65+UQSU\N1-0H\Z;cF9>I[X;WcfFU8U>Le7&=0]g_gBRS=-,PecP60K
cZ>@EG+6:J,8&K.)Z;4L&P<-9aKgMWE6PZ@#C(0PH)Ta+:CD1IRE8&GC(9LJVG]N
dA,6_N>&[BecY\#.@\9P(\R<HIXUdAJ<>8RM@MVN?ZKbYJY]6(6+6f(.DX-/dZ2B
?Nb3CWSDcJO#Z4[\AG4P2(,K[R2?YA<Y1>Vb7,ZLAd)?-X9.&9DgY.aVZ.GbT)^]
F57:E\:P#QUX5KL@eeYODCHWM>-<=>5a,G=(7gQJ=a8=I@PC>,5BE^,f1;gO9?H0
#M[AC5a:Xgg;SFEEW_dL3U<af.3Q)3;#JWJ]aVYD0_3-c8#5,,[U/E5d:WMg(bX>
5KE0?XE^TG_)5cF1-P[f><0BK\dP:dL/T,+91:FaO@&F-\QCeR:/7PC09Y(XP+\5
VYQ[^?NBTG]E)YP-e[P+;g#V,O4c4:I)>2a[[[.#MS];,eWKdYgW_.#b45fGD3<g
MPLK5?A/?[-[4E,<<_/gO[9(,\UH9+?2c5)cfM-7,@@\H;[<EJW#_;8GNYZ:.F[g
V/DKF?;0I_?d(M_U:e:1[X>CVZ=PJD;dD?b:FdKb,.[NXM#U#.gAUdc--b,[YZX8
L=B#^Y<4=a?YP8;LKV408Cd41/E,XL2,e5K?#aXYVL[1Z<#C98fN6+f1U<LbJEDg
8(g(X=N4?5F<)Q69PQESA?+cLN4R+WX:,-.PgaH\\;G;&(5Q18;7&R0_=8X>B\YM
[[>M2=eU)_e,RS=]1/THKLJ]MATF&c_=4K]Y#?,J=16YK<FHXGG<VR)4Y2#X_CY?
FZ7:B\HTPY^43+M@d+8=YC>-2&c^19ZY4ES)2YI_;dbRcLPDg3dV2Rcg?&WB9HA7
.T_ZdJg\6I?_D+P7+.O5-U#.Z[7O<gcE?/QcRNR:@:6O7RXF47;6dG?fOcRSU[(V
0d.2X9f9N.Z^&V#5ZXe1dKH4a<X.:B[;9g+JU).-)P?RVBG)RBY9.8N6_ZIMK9L#
2ES:gY(&cD,f4)[@&c,0V^E#NHKF)<<,2<SWg2>Hb]<6#^\(^O+NbEFAI>X7TDRc
W=D&U=^fAI5:1=_F(OT9.CQ>YDI2UF_7\]VJ^P5&(.KKQ8Q<4]cc@d)\SCW\b3?\
7XH15@0WEX_AYd#LaN7aN=0<G=V&V6(TUX(0;f^SU)J,2S_V\+L2K\C[VTO(TI.-
:b#e3(\V>J.bS)^/F;<-bg.84[4T01^L(fc8(4@Ab:8R2&;WW9C]0&b6\9+H+GR2
OXS&g<\^QH68)0/.[?Y30^Z@aWXV34gK/.OC8L]SX.F#2\-0^P/bD,>Y>NVPC(OX
NE-V78-IR,W:1LO+VT/@#HCGWLfOg\+B7N5(<RLLJO=+5[D/I:]1-gQA4TTP03gL
;4XRZ^A,\O/(^?4g=:URLQ71Ie]QT,+^>:SY=4[+b1TdOE9N.)+0:-#YdO<P5O[7
+G(GcK^B.QZE6KYc72e7>.M:QEKXCVAXeb9[eAFb:2;XF8<M4Q[(c3cL7D/3ceWZ
WGL,\E6#D_.XXH4Y;,T4T<He52)9EILTMPBg[N7Y;02Z=7e&H3MH(LHZE&(ac3_?
U\^#0UHaR6?Q3;@AM/:<XF.&]Tg9+:a+(eG@eeYOF14@/^NJG0+6Q4_M8&6,-d;c
-8LZ=CQRSCR@3e9K3d95GA>8De]9fgD9Y.H\+Rg0VWO.K:&Q?X4X9\91MJbY&O,F
[J-W^_B7,_eOT4(5GbL^)bQ3c2P^g-X[IEK/-?cF1&DG3=0EG?^TOg@=:4LRY.Q-
QX/A?<c;&+@A(^0PAL.V<UfSDKWN&HTCNA54C8BGF6B0e;2]eabAB#4\[M/dSaYe
D4&UR#5W^KbFc)V3R4.=DYFSEM01e=A05#?V88]Y2/UR8R:?3HPd\_A,FE3O3,FU
@NJ^)eAf?R>g;fZH+[<ScB0J-6gc]<8L7>F?AM)JT?cRCVFT6gLfM+H/fR.0FB/O
ebHPOa5SZJ20W43(8g&>FageM]2R+?ZLDF#6R)f=^,9Zb.6]A;QS,C[E)B1<aSJQ
UDLF:1U>+gU?E)L79+R64:P\[f7IGTWN:#PT5#1>fVeXO/V,;6(9@0MC?Q>)Z8Y\
+KF=Sc.XfFX5)V;+]4NYQfJ2-9>Z?@Z.9&50A@0^,b]g<:gJ=Fbd&dd<;FKaG?DJ
=NMA,2D[ag,gJBf+V/D<[>5UAB=c;.\XEbDD0VYD+CCNR&baC@Y0FN:1T>E&2(g5
c28)U<+EE0g21UQINK.8aB8I48/1]V>@Ia;M(5V-:)&[ET6Hf]5AL:RM/:D9f2@I
.@8XH^BV,dFa/Y,f88Y?c;FMG9+/B(IC6(R7HD0QTe(_]UHPN>fDTPgV&SK_JRY4
93;b<+-:,;V(HJP^UGR&F_D;9X)S1cYc9:KV?@+c2QNM(b5?:<2@=ES0>Yf)J)#<
:+R9UI5J3faZB=(6C[(gE32@@8],fbf2e:]PHLP304MPWR[[XCNNCWSLc9=0CEaa
I-+&aeMTA(+&/Y_?PN4</F\X#cGFe\KgOI/B:B=J[-WAHKL/U2&JVN2G__=5UbE8
G]7aDK&b[e#(Zagf]6:]S@4?;eZX,Z\8ecB)Q4BM(5YAW#8H-[92,M,;PDBg^#B3
KT8O1(VBJOTU0V[H9&F64:g\Wc8#=R;^<6VPS5ULeLZAJN]0a-K@=aP9(]4X9FYE
88^d)TNOf)C3[YB;ZK.HZ\HC7=O6OP]3PN5#a#-:DP@/J#V^+_IOIL[#f4U\BVQ@
EWgN/P<Ddf^P>V_X<E9\QKL+R/aIc8#3(6:^J:FBJ>DX49;E&)7HFI]JA9a]XU]A
PTcgd+YR7YJSQGZPZQ::&<V=>:Ic,3M6f4H(-(/EQN\.B&FHCAC_c/J<b_P>eF42
W2POJ[5e>UdRdUIb#XZ7XW76ZO#I:73WB2Aedc0,LT+V&?;b&@>JNQT_]g.M1<Pb
^LIMdeXREL&PZ2=O.]N3-7_UVL;c:R8[_TFE^8(]+N2MV))Ja1KNTW?cg<W)<U&5
;SRYRS/(L4)O[a3+/N@#:W?9gLX(_CPB(LG]Yg&N(<SZM,&ab2_83SH/A_+K,bRR
.35V<3,CW3(B8X:CJ:a.X:QfB),McXKBQ/NXc6.\?L;E;&)E;PPW:BP\?aZK,V;3
,5X[,2GMNS=([B>>Q1#OKE2Hc?Te9<2NZ01Yb]MU=8YL0)Y];@LF0A:GH:f>SbZ)
6-7V.-4&MNTK)6P:)?0Jda:D9ZE8#97,YE=6K8Q+3>1@WEU=<SVL[@5c=_f0ebQR
E/cc<0&1[g]DdDZ,H1Uega1HfTXNMRg95dHMEfEZ4NfMdH<J)gAVS4Fg=P.gV#SQ
/0T,OcaK.4@2P_1WWF8&\)9]HXD>9KK@0Z1F67_9,K5RX[LS:KD4-=6\>WTW4MS6
O&;P/BD:MPg3bgeM[Lc.&=-g<cNF1+?Q4X.aG++UUMH<e;-dRH?-4--CWaT1J<@#
:<^1Z#/7S,O9bgAFY:JVg._LY8RVQbWYQP#X)L44&>(,R3_W6gU@O<\8Jd^a=Wf=
F2)Ke0;+;a9JDI0:3I7CHAf/H_)3NU(U8?-AXb#R1+YOG\V5LcF,2NYML1D>,62K
0V&LO([A;##:2HE#JH63dI.>e;d]UOJW7Kg+P+_e-BKUDbKC.a=)KGU?Z.6NDZGd
LV4C6->\bXNQXW^/84g\&GETSFYB=OZ?IRY4NM1f0Wb4134cM;N=289CHNF7CdKA
CULbGV9A+ZZG7cMY2^#-)7(f+0RcQ?WM[E,E.]3a+gGb@c8Jb>X4b)VVLH.^:8[#
HU9L9:J6b)4AP<[+We,GNF#ReU+DT.2F;a4\]RAUZTTS/HK@/8ZIU=b#MgedUc[)
33/:4N.^A.]Y?)8-])2/IP(a8[6aeIfI@/A^[<XEPD]I3c?I\/.ga-,ES;E/XKg.
bT;96(]6AWT\[X@YP05CV+#8NZdZMKLMZf\38gN.#I+EfGMV.7MfK?QcHBU&>2F#
b_PA>U8BZ;M153HE.D2U_?CN&Q.2XfAg69c5beRKM,Ic^5,<R+=?;.b]<b#?:A?b
(K#6B@KWP<f])Pd/d[5UK,KaW]^G-)PNOP9b=5cfWBUBJZ/06=D)?G#^;&+9Z:/L
P<Q:=QXNO@d0gfT:7+<DHdVDH]/ONQWY,^X.6?b3Kg]T7TVe628OAM>3T@#5NV>;
RHB0N;#RT7/>Eg\Q5c9E&^BESAe\V\4^HWVB;gTT@d\@>J6T63UfLd+OI:1@F@6G
BF:Y\3RCgUC7,)33NR_7(9?O7U;\dJ7YX5\dUY7XH^LYD04=W^1K-W/,eY-,A<H>
=0[-(J-fLcG@FWJCX6<U+XKT:TMG<SUM<Ra6d]fEQVFYV\)9;Abd/.Z+T8GOLWG>
U2\P;)JZ#<GP]I=5fRI&Xf7B:;0.CfBA&<@KC9WELEQ>3S9N0c_PTM860_&K;1\L
U<VQIg9>GeN()c?B4E8TDS#,Z4S(NXO5,:^&Q4I>e:GbHT:\LG]4S)^_.75YHX]d
Y5J44dEX<,>c:L]TaZ3K:>(6ZaQN-8.18GZd04(U>MJPYLWRbJ8;&IL9DEL\a[@W
[Q,Yd/gOS3fV\55[>C(.(AaSbJIMFJca]^@HD-WW[b:c6F]WBGRTEE&.,L75Y7OS
-;OP-d@PMF7R[(K:cNH:C?EP5FNS6^,Qc5?,#=7C[P^(;g,g_G^LCO,U&aSI:0#6
Q:b/)H=@@6)(9S=/Ra#KJ6ALQ416e[[3HCC1-SE1.2c()PWT1N?(2ee?KaQV8GV@
Q.AQ<a3cbeMMg(\.=GDC[X3:DE(57VCf#V>baMGW62YL:(9N333H,#f<6OH9#4Ba
C\89I@)HS6CSGK2+U+]b&c1cIA-.KaKeR.:#)=SOa0\Me\dZ8FZLKg1FHbe<+/H8
L9/eH\=Jb/cZG?GN^RKc2Ie>UY76>&^5ROZBa5M44N,JS>4_XQ]9=GO7&&fa?7I6
VdRMKHGHcKC8#cgG7_@YT#\AA)7U:^N&0TD)1E_E8bbE.0MeDEITF<>TJG+<H61Z
X:]Q/M>)6JPIN3d0YUVMY;GQW<P@LBTO(),W;SUaBI>I1\1AC)KZ_GQA)=deKUW#
XW=&&eBSYZXdIDKP=(L#E/SEZgXW[Y_#YT]S@I9\_6?Ve>9X[7Z6\99CC328dPO_
+OJLWZgTcLO_b4C&&Y^N<@OccYTO^J6=dfI];A;3OLGL-fZ6T/d(.>:)bVVG@KGC
S4]P.7H3T^_X:)d&eZb7Gd=(97\2adMN6T^B2:\36<;JOa5baM((A5fV:\6c^&HT
,WLI+8BHWA1,)]E;[0ce6bb4OWe#>H5B[ZFG(+26TNZFFRa8H@:ZL.@CO/:E/1(@
1FHH9>#SNFIJf.ZO026]JA>@g[X@FeJ2]NBK6EZU);U)[<73=-WEHGO<>gOZ2@QM
??^?@/6EPb=KQZa?JCO3SO\9?AES)Yf,X8S4g/GD1\e6W.f-R]@-eg)f>MdKdP,8
12)KDJc)4W3^Q;DA#Va6?+?U.c=\7R[PU_,4#W^<.<3NER;I>DHKP,4<KMFLdBSf
S9\^GfQC=:CR-=O&2IWMTZ@@0]c\\414=f47bTU-dC+4<9BYZ#-F=Z;K4GN9&7(7
.WHVaP<Re1_Y6TcN5ZNCd+?EBb;B6UYfT.,&[,6BaSP<5)^cLb54+>9C2<EVd>J)
-e7IG1JTW0b=W:1Cg-P+LM\CZ4V]8dIY4J6a-Z9V.Q/_5,f-BYF,9#F<ceEM/OJF
DFba4=7]e:>MGeeTS@R2.8J6(Jb9WC;<RC[D0FBc<I(^=c(PaXR6>X[MI+?3/=KW
P+S[7O1c>e9(4=D+JKQX[N>A4_\)GFYEZP]:5G&\V=#DIZ])I_OZ+Q-c<8:Q^IT&
3T=DQ0Z0MI1DNQES\O32R,3V>U3K:EHId)XWT.9Uc32D@Xc24(HB4W#C?&VWfVZX
N^gC2.=\HaJdR_Y0fK.g/[=+-+&XfA)5_K?X4;ba<(Q]+MPP@C??HN=UO/Wa=e;P
Te/HW@SgaLTO9R)Wf2@Oag32_3\9\\X:&O0SGF\aF?WS\Y[6_<Ze?:+D(fd(:Fa?
RKC7gWZ(P5]Dd1=#Xc(1dMK_\bHC7d<D^6^L>VB?,IZ.P6d,V5WX&G@gDOO6//g7
M+#B?eXNW/HAG9>M2gU;@a=^]ST4@TPLRZ(#K^2OQgbZD,Ee]]_P/(])]+.cQUGS
?cS#S)YYIXC5]3Z=CD;OEPAK92dWY;^Y-fP^#YS]eMd)5TeeaF/&Jc,(BY2QaS](
1N7K9<KEYgcV]H:CV0B.]0g;3(0:+7=2MeU;/#?eM<14GE(U7B,Sa0:Hf)OW5U83
BYbHJ#gIKUYZ^fd;Z67>Z<\#;71?gQMe1EgJ1C<0D.B^aI<d7.Og)JLM67F]#e[3
O5)TFc&V01He[M:VRX_E)&-C7#6/A/>H^0K[PP=eJE8B9VDKK/M-IcB@@OA]55[L
=YPU(N+C4-E-O+]T(\a2TZ:?M)=T)MRf<ZT_8D##9>]a[K1CU->U;&aTXb/b<@LX
4JT48PgK/CE,R_BB3G11]N3]TRE6Cc.)?DM&(;1aEYAGU,/,D^D^gDcDM08YMCL,
-/]HC7BY6bc-UF4B6L\Bf=\N]WU@-7,aY5GN7P[RV?JU2X;E-8:_]Ie/2;+-ZKU+
+,aR6faf9.9PQg3Pb9d-12(b2N8fJNd0N(cNL-X4/_##595:>MMbQ1J\7-PU8-Z]
)6_BO7)>Z:3c4]DOLZ^X;N2L+^-Mf\0_D1(eK<_^_HdFc._0=4\MC]UXFIDWaYLD
6(P-Q6R>J,gO_B[/WNEXJc3?_.?PWW=[389fZ32<)OM>7aQcA9->=aUFb)9FDNK\
B[;(OX@9TcU8U14Z+4GefZ37^R=1b.=OMa02N6fVdZ14ceg=?YS9)&VOUPPD+YC(
6aR>@>Y8-)1I)C-M;-ga^X0V[IN9J<>(Cb4;&,L6F,RWPSUc(X&_+KL:bO.eRB?6
PZB_K@\+>)&f)CZGMd2)GH23fNDg5,bef3<NgG9##U>&R:PPT9X1A)QXL&+;WTIP
CFJNdP.gFZ,U?9e@DceFGBSA8I@.G/cBXN,>GG>@FM>X/R+c+>P3):7^?:-[MaaV
0U._P;Fc>/I20.H=UHfF,_XNBG.:3176/55;^Beb6BQ\_@Y-dB)C4KGV@Rdf&U)V
-K8Pf):X,Z2DQafCRbf7[F8^@FW^\>YZ9YbbRb4((a516Ce@??OabLVH.a1/RbF@
[4fYa:Q(#\._gQR[J;&CYCWFYP@?eH(/a2U1KJ\dBcDEgTG<FW,#,\M]_gQ_P.Ge
T@F&[d0cV6-0AYJSPH3OFdNg(66X3+GAEg4c9-bbQP(E43[-@RS(^DY\>e3NM#]/
P_I+@H?);9:0L81)Q,:G>]U12;Q^3I8NQ^NXMcR12=>QN)S@[d7f4J[EVD[FR=51
:3\#aA8R6WJ^RG6SOY)Q4GAZD,6MU0CdJ?>SJNRK?A^a;KMb+P5Za+)U_TC.&U5M
VJ3_AU291^^cIEKJT+dVa^:]A0F\;4ED)R=GE[CgT@44M7V\9[A@7GS?Ee;>/gWW
G5D4EUE[0J4HS;KR>4^9f>,YbV6Cf4RB,Ie5g[B2EPJfWDO>?&b,F45W&V\W5V=g
./=+=X(,^77f&L]I<4LV3U@Fb#TE[Q/DfLVCRC0CG1IMW]UWP4OgRSC=1(e8]S3F
H7gQFVU<YgECL&RI/QB+E.^0.<S<7.).a7f^544;EWK:RSH9G,3P;QDN_A[ZM^Ne
G]3eM:T4@^Wg#GJgMFHX>UWc@fG6@bPEWd=7FFaRf54UQ=8.dW,S_2CCgLZ]UHUX
d)aEG3D/I9:8fRPNKO[aL#Kb<]cf0;K2abF+:UJ1F#G8\e,^LK3VWG6\-@EU@-=R
W\16Xd;#QMQ7_T[#650&UE<+6SWDT?F-KYSQa=-9<&_KgCS9;f:WDVQL4CECfB)D
8><b6)K8BO)1+BG/#0]2fF:E=DM(T)NY+CAZ>P2XP?B>M3&JK/)AP7?aTN;[DJZS
VZbVT.OA^S?&)_0,5)M..+K/BE98#>\O]+0MC-./7V1\cP?2XX<N5FU;#@b6L(Of
0./Qc.94Hdg.D+(?[0UU7H_a2.Mf383G]:R=W?Z)Z-)?6\]R0JSQfeac=K?4^f<V
?SLFY7?2Z)1Y6D(Y<QS=)1>1B/+<gc4cDYK0?]7gF55JfL.N1EAg&,?C7:F[-aa@
7^INd)Z_B3JEB:UR]W[NO(,^T<Z2G;G1<P:MY7fAcQA]OGNEP7fJ,d?/Sd9)@4DS
#CWHUGDALT1Eb/2LN\9#WEU\=V7UZJPcc6/A;g9JdgT43C1CU[T:\3)DJ?Z._f][
K_1<C__GG##;)J<W\RZT@M9-d5&?e&&17Se>/U?TU;H.[6@YN0O>N24]gZL3<B/f
#3/bXLA?U]KG1Pb.-UMYe:1G[8BZZPX<<:aY=9VAbGaYEV0W^H;)=F@dF7XSR:GE
C701+;&^)SYH3bJ56\N/HN71U]-:.Wf?Sf?.&L5RBgLQ>)b_0KD61-67d\#N[NVE
.eWDGN+34DJ8QF_2QW[=]Xc/R&OTDS6,T5a>O9&L.)e8<P+RO(.E,eG?-O\+HgEb
=_?GF/8P\=(>Z-K\2]S5J?=(?>68M,7HT+B#YY@<<;H6=&aKLI/b15;Y)2LYbNZ6
Y+KS+)N_Nff-^f(;2L6\B.(Q9TL>dacdL>9cLLIB^QK1<-,0\#9CZ2?Z0I>FK\AM
DZZ?[L5-PVV?I-^TULB?6PVH@R\J:ceR4FQe)PYOgIYU1MS]ba0SH\D)]D?P@L=g
(Aa_4=?6]2db:ZggV:2GYPgM:[W^RJ-9Z:cbNU1ac:-=fN4Y>8^]]:[>;39eF-=+
X#QSfST0U,ef+GHE+3+V>A28S]<4BN4]OJ=W7Sg/)X#c,a?_d(@C#&?XDV\cZ>W_
7\.C&61d5?K3\DP2V/F0O<#\feLea^V>;0O:UO2)OI]47],MVWb>HU<_,\SUJ,<P
H^E;)ZOdeVI/=LBM^FOO=?/(3)YO_V-GVXV,7Zf.@_/>4@P,P&De?^d4YHQ>L6Ee
?YgTR>M3SET_dFIT3)/cLe(01TVUGLaKGP8^\Aa2__^_3dL]A/:EE&gWE0KJYH6/
<+\g\F[CMa#F2H4DCO74.UITSKd;7WHddB/5_EV+-<d?HZFX<c^C0#.]>HRK=ZX;
/16\N=L@C;2a]#C9e]Af[U9L<PD4#e^9Pd6FHI9C/&7BTJQ&E\(Jf?[4PR)O76X,
#>]3B@=HF[+M9aOHA+U\,I8eC>=LIHWJ89M46>F(=JaG9Q9P4@=C&YY&aP/=1BV[
4@B#7=-P\4b;O0OHgD^XaGXWPPFgMdCI+&SeOHOPb/UY8[T+)FB8MgFG/4G)F@;J
I]U@R.VBLP-f:HK64)-egQG2I6P(#A-=3?2ea<2+^YE12Od)G=4JIZ\B5,LO.S8F
T),-A[/_F?I,;W8HR:C9.WZNFRB/X?>R=_S5SbWTUON_CEKaH9fXN?#a/O;3F#OS
?BI.XT,H#1>.O_.I^2Dec<3fJA._ZCWVY9b-7&-_0bG[^V@[1[T@;6R/U;M3TTSY
cNE/>fUC#HNe1RT@(=Ue4TR/Q;OZCS/[<K_)18g--PZ(e]4;WXZ-K//abJ[3228E
/F7B+X:<Fe0_?U()I@6:Q#C-_K/(E0RaVT^J,ab.gFfFYgcc6I#XJcOVW,De:a&K
#O@[0dR/J,W05^09/Oea5S^^<dP64dH>Q0.Z,NA<VGaO>Ze-YND0T.Tc<7W&]6BB
U8b=X5\N1Ed3#.JE:K+LL0K,(0]Z.a]LT5ZA\gW&^9DB)2eRY<S6+#T)>I\Z_NYb
HfWQL6,(\4&>KGKLZEB5WMSIeG0UM,ZS)VQO3&eT)DOW<4WPT+ca:>8fIL8SJLZZ
JX)VeaOXAD>\Y\Y.VMZ\BIU,LK5/1e+#;T3DD6g)@Y,&V[R(eL\Y:M7))]+<Z>MG
9d\^V<6N(&U(O?Y]OJ,7)gF,YVW)CRc&Xe>=>WbO:Y)Ffe/X.&eUB;5/EJ(c#RYU
K)??OZC06B-g+Ed(bcG9fSCT-=[\>VEK44F<C&gDVQ[3>bYM[VLD&<#;b]cA@d0M
[aO?cBa2?Xaf>?RUWU&0A=7;eO@(3&b9XfI)S&SU3.GcedV[IRYM4N9)c40H2Ve6
fMIg+..S=WWJHK4B=MFGbESb0@WJMC2R?b(e)G/DC(aW)/M;bY),f_3PU:7NVHdU
)VHgGD]@X5KWHK+FEX^.UBF5AAZ0b/U#.KN&B#B4Gc4.=_(d==Z@TY9Qf.)KG]&7
AdU)G>-<L4^L&63bF:W<1#-CCD&O<WGc+@-Z\FEY;+@PE&Ee><ECM<;FJYY5@V3Q
c&-TeM?d>KS:N]NJ8+PdUCa9(f[#eTS[eW]\DM<a610_R=+<F4d3.038NJ>Od3J2
RM;\2BM8IBQ[#6WJe@?V)PR3^fO/R2LVOY@g.BRR@2[),PSgP;89[G[<cBBbGZ.b
(S=dRYPR=[H?bVb1/6N.A+8C?0RU/]@HE_Z:;WaGU1;&PX5Y13H<ZA?TA9EcN#Lf
G5BX0(?/SCTN_a]LY#5b0;;e;gF^C>:_dV8+[J<;4L4B\X^OKb0_X,,I^dBU7d&R
^=N/C;TKXJJRSc:EXEMIaW]D_XG:A#Y+/)RY@37G^S7I.Rd2T/_g@b_Ee;)M4^Sg
((I4-Y=4#Ng4HKV+HWNcLF7b>D\b/=]A&,EW,]G,J9H-;;:bR)SE0R>Z>gFDOgMI
JCHe&2(DH+PU^7IK01>b,KIY;#L__)KG>UNVKTF<CVQ+d-/O)fCQ^K[@e;,c7TWP
eZeeLTO@7@\Q@#O@HPY<]Y=M](Ya4WC63G7Z&5V71M9.LAf\[J:^A872d+9B1K8X
2f?g7Yb0;d^C3LZGG_S:ISZ>7<EKID(E#D2F#ec)BD/_\N7]e/@8cWZ-L(I>@22U
8DTcNZ__3]>?b_W?UK/_9<]FKRI4eZ_J^/Y5ZQ+)O4dNQ4APVgX1&g>R]Mc-aHf.
[/)XIc;0>F5^18Pc^^3Q&KeE-VO,@d.MAO(YVXHP@3g:gd=?Ve4S\&G6;PQ9PFJ\
fUd7F/NQ4SB;H\SWeTHLEHJUeWc-ODed<LC^4HIH/^a.D#X>J=<WKICNR1,BdPc_
^<=Ub-:WN)^1\?3HVC_<KLH^IB@<5gU,-P8[AVVGVRGUTf@Q43EdX;O8>Z@3FD=(
0]J>>#6_Y4ZWege6&&9Fff1dd+aQ/0)Vc4=DN\g2L+cA:a8g&3/g=f=P+WUe3a\9
f;;UcH\;HXEUdE;/],bCEQTPe7VT(_^+JXX0++^;0&F8G0MHG]CSY]#Gc?=//3E#
g#Yd^W/e:G?NMRI\M/V9<_T5@(A,eO4/>?+Z?9L?LdOM<d@]a>?M-/5<FFB:-QGg
&TO=VNa2NZKBMWE19/M7=7IR0&WQeJd&e;33a=.?G26Z2QL0:g/X_;0VbV:>66_D
g73W+M4,c3+26(3\R3V<[>f9TO89aK\9V3Te4-gLH9_U&AMC=?7)T^]1&-dI-KKI
E=aYc@Z,GUb.Y6/]^BBA#a2NCQ<EJVU]g+^T:MVF2GTcN(6gQ.>/B2faNcQ.X[?>
^S48MT2^DNB[ZF2\?_8/:/]D+.3ea=L7FFSE>,\]6FX:)W7)B-3;<^bM\LPaM.^J
.7+cPARN13Xf:2V.VgHJ+dH#Ffg/YL2;<c^)BF=&AgCIa7M)g=<efNX;VdRVLaB6
+Baec^#\=O(D_.BS:BRE)>)^0f9e,?4(PQdU()?(90AV2FM8d/2[#U,BeNY94a0I
O53;?.VSZ:--^#(L>aUXH\5H6A=0MI[8dDd9)RWM2H=_d,W^73^.2Q;Z_?@LV,bV
]R4TSSU,g^g3<W@XM(Wa-?;0/7/,bgBX[]<-FAL@O2XCI]Bb2O0#D:RB/ZG#f3:a
1(18^.4U(0BID^O=^>X9Pa60PQA]FN.CF:41&UH\H[RG#2W6]^U:Pa0VWU30+^^K
QICc^PWV5d\CWT0>dZLL<Uf)S;<HV_?D[(QgbFDM9_a4IHBEI0<_I<3)4f)Wg?3Q
#PQf+TG(QCIO:GQP2.g;F@dT5\KaZE>@VH,\Y#LA(VWB(3EHDD+5WA;D?B-J#5/(
0=0Ae?DHe67RU?#MWa,eYGT:&=7C5>9-C93IHTBDQ#XOK#fZT(Q3H;8G;Xf.0J<X
[W,4f^?I8LS3:8V0[;GM>Cf7)##7+:4EKTe5ZBZ,ZI#JCb]_^IG(9@I_g_P+YDB3
/AF(LIKCAZ9[W+f.BL8W:aI];MLE?KG0@WB\-c.G:=UP4J)O:d1^@((1(DJ,\f:g
8J&)M02FG&)^]gVNafeXAf^Be@=/0(J.8;SG^__@A:OM7Q2INBNU6_N2C:e/^>XD
Y&)NcVd:12P,.c-_JV6dK_)GSPN-HFeU)_MSX-E,Y:O0YR+]&>d&9McZF,C@H^)[
?aK[X]>BFO=\4+<,;T9@6.MMgAfE202^2Y=9GXT&K,HVODKGbWGA8WR1VYVT.[bS
;(?U@C=eW.#66NL-fM+MgALeV?=ge0W]#AEOSN57PXT;JbJ0N;(1Y:VNGJb9?VC,
BQN6UR[TWZJ2.9g0C9Y\T_/(#Eg923#F.U:NJWZ[;H\]))I68^VMJH<@_:I2UM+E
f0<2[=Y_=eOS5X/WB4dS6\\<<b[UO@ECe)25=aaU)S^]?U10.3?:1KPB@?.Lf;X>
&aaN\7[28#1S=cb-OecV]3]gIFO/+#)Y?a-+C\A=C-TdA-,#)f@eQCg/3):W-Ha\
Q+H-g7gT0edc3]bKVSU1\.(1_;OcWNER4F<Z_XbIg1Jafc7R3&FSMD8@<^B;Y/,a
TP8F2Y8H_@+/:75WZ[1C4?^Q3ef7eO>g-.7M3M;,X,J))6M.,7DY,Qfb+S,\gIL2
ZRMf<&R24U).5(;O+CJ-.&JRL(cA:aGE.E?/R(>T3TGg^>USbD.^^KGVM2\Zcba3
FLRAWdQY,Na^e8:^e_T=;Z_7Jb#L0=e(=(\DgP,2H=6=HI?DK)>A\<..:VW>57XM
Q[0/R]A3=D#QUK:c3Y7XU]RC3CfGIQ:Y;X@8K=b2^+C/5]<GNeGL><1WRRN\TL,;
,?5:C393L>defd(O&)9K<R0DUT7Y-?+5c4C3LM:VL4.U<+)d+V7H;INNBMgNIT,I
8R]J/V-eWSG871U=;X.1SY/fH-;.Fg#Q[#YLd8R9Q>0V&)SQS@,B\L-.6Q;-8O(T
.POP3HLXRc&M1)e=CNPL[+:<b#R1([d^TY@T]6]9b3c3[/A6Xa>6D<],<Rf77F5>
<O::YL-1O]e;A9NS6,;;2D0IY<8B-,]MBIL-11:0845MXASUf+KggUWX.0/Ed&b5
E0HPREBY1Yg0Q3,@?2VB=)g[+7,H;=I:e6D)a.dX5-1O?WHZ<(K9N/-Q:aTX4AQ]
RN9bHc&-924N#Ic&Pd8RZD@7=2WgK0/;K[c.OWNS/:_D(-1:S?_eZE]<d)(fX4WF
J,9YZPHM=G>bgd;IZRZY6+YS=G-KAG=UNf7:R>YO@RL\N,]:>3CA>f/3+571d]\>
:>.F+.b>B[FEa1OS::Sd#V-6=R=TI]&DU6]73,<NQQI,07&VFF]eFWZT4GV)W@J\
-XdMVKZ.8bTegQeIB^,MgCeWTBKcP#]WK^QO3Jf.:#,&(>BYOE#@E/CBD:;f?JM;
MLJK<&OAE#,,E[MTCc3M7.9E.<7J67AK;7H;-:9G:GKc:I/A8]c0?KY][BeVI,-X
]?.ES2(WFF&E^#ZQ:NDM/S[OaL9B0->(JP.=g-4F1:eWQM<[8_@7K/NMFROXdX98
fQZY.2XUC1Q&;7fXE0C3C)A+,=;7?-+Y->Pcb2FJO@AHX6Wc-RgIP#X+WK>GWC3-
1BN31A\\HdF]5C:_#O5C;=T_?>I@dLG0>+7+O^BII:M,+^?aL@DK18+U<7_<1Sc<
/-<8+H,N)<;7R>]T,UgCRHK]@>-b?.Q97@H[1#a=/)8XW4MMf^@c1^3\9_Gc2f-A
N=DCcK4H>ER4-+\^=)BVC_&DZYD9Pg(6MAZRP^8H<KU]--=0&H,@=d=K4=WZJ4.0
/\DW>BdF2?g9_[R_B&JGXV3)L_g;fZA#f^/Q6?LGR53Q(BS?FP;0=+<^,Y(0X#5Q
/c:3@C1@;&a3Pb?&Ye=-6\PG^3cH;M5IDLY:)?cGC,.<;IYVIg7G53V(>.>3a+@[
A\T]A:S-dXQG3YLU+05Zcd_Q,>=P2Y]Z&L0ZSJ(1L/A^.VAccPA,X77_I,^9)_f@
?Fd<PYBDSbA\C/8Y>)Z;C<ECO<6206R,E&]YT;B?U_00E=6L>?-f>6CUCQ#bGYXU
GeOEba,?015e&BK2H@aF)0[(G-4D2=gb<eDMb684EC#;8:6/?]bg#9R^-5D1P[Y]
NJK>#CN?:(5MHT:>AP;G:0>W,1L_6b=7CS,ORLA58b<e[D15F-UD4D)]R@6LK+c0
^f/FQ81JJ/:0EJIM7aJPA55P6V]XY9d=2C2NT2V#C0\QVB3OeXd_-))]g?KHb(R8
<PdcGYPNAM,J3\8K73,P,3cR5<JcK\T?A99;fN\Hc&CB&VGSRN:Z_1QV1-/VF=eN
XF0;G)8)\/BU-R;8E.a[^73,Yc<JNIY^:T^YMO5MeSH0]e<U)cPSb@A6I_2)PO1f
2>+F[&;R5M:4482b+6N7:2Og>I7\8A]U(J>YId-(b6/DDQP4@6=734)4HDV0T]Nb
9MEH+3;aAS-Wg8_H5O,Q/2,[_,/:C_NB8KMM?<Y]MM?XLOMbI4T(+[=EDQUV<(GZ
[2]\.<1?E@R4<N&:;5\ND3ZS#BU;IRZPfa-OeS51&Rec7>R\V/NNI81/)Y/^Z?\S
^]d=d>a#,f(JD8f5IEB##0=EZ=4.A5XSR[@6eP+\0W5g=gARg#e4T@,O3WLO=DB\
9K_8:@YU:<[<UN(&=6VWX_I_ZF:YCJV:>4F)H8X6bc2S)f(Rc3(eE^P/23)8F1Y7
.N_+Y(DNASQ3d<X0NTC<^S5>\B+,V-EAG)@Q/TR@GG=<K3L?M>IU8bFEc\AW)9MZ
Bd9cR[(S4D]PB[6JZ\EAJ:d^KQ#C,@Z3>T@&\L8S?KE2:d1K?cISG;LDg86UOD\L
Z8]4X4N=D)[,CgDF\OFU\NAURP&4XNfSHR;V?R^Bc_3[CVS.f#K(4M2[@:#)Q(>9
6EHbb2,Q,V@eA\PLMK+2(0c4P,W#16_3:K@D1A8dVR;H,T&0BSTT\FJXBVK.F,5S
3[T^-X0#.N,,g7+TWe3OEWC37<_UKKR/N5@Q+0([U^EdU7#(abd(ZVdNL^#)./3\
5VfZc0_DOacTB0-g:5>M3QUA\[?&^S1TcEI^/EI^=79[W1aZ+g(7#DX\/^bF75Pg
/c65.4@;REEK5?JQ<Jg/7V+eH(#L3B]7UBJGI)IO8>8^V7H#Q,+KXQaD\#586==B
=,=b^47EE]+0_O9=WU>RBB)McBEANDdVERVNF&AdO5NSDZIJ<O?+TbS>c&N-f8-+
[9c[f9aEXAZ#JGNHMGT&aL_bI1\DL8g_X4A_f8#<>(e/1C?<(GYA<&1R._VWKTZW
C94Q4+D1b/W]8B.Y.D9bL/3F@CgV/gQ:cd>U3T-7<.7<WNgG.@ZP\4.eCK:bSFMW
^E[/R/6BI#^=S4WG]gCe3(H4Q1>DVaB/W8XN=Z-ZU#E=.gF,H;G4XKNe4O/](0AZ
gO:\@f\]0f28&3J4:^>&X?e>c&Wd@[[d(?f1&BLJ52BGQHe;RL3>,RSOfHQe.O6,
^FO,OX+YBF##;=&&^RLZ>]3gCJV<[.RgS44EZ8SPJ>C@Hd[NO(YI_BXe(>TO>BcM
K0XH\>OcPSgJ@\IN(.>1&IM@OC8_(:R0+K]UZYd/89W-N)9H=XR+/U>DLcE7DL7R
7Y#>IfN[SfY-UHF#;TDNFVL-?_GR:cN^aWWXB.;;+N3>J(Y]UHKRHL,CBE>NK/>#
g.[VXJfX_3@Lcc9<7T/9Q0T7d2JD=0Z?M\L?-ag#/KK,MU_;NdNLH>@O>LV]>3QB
6Y,,f-ZSS@9:;(=@NVP;/?J-Z1U\>6S#\[e&;Jg+:;-AI=./4@;^Z]W6P3385O_O
;ZHe2P_GQA\7bTC7JHDE8E.2JJSF#F6APWYU0AdH,AeSJK-@D#gQ=@3UK0V0[;(_
2E.cQ.5fUL:/)0W[1C_M1EB91fZ5YD(Q++Y?.@L;[6AASMTF7dYV7M6R4X6(:eI0
CA3f@_e:ceKL6,H5@fCI0D6Q>9G+<aaS7[_W(86c?[OAc(W\X-W:U,I48R=U?U(\
,?)D?KX_1aU^DJg5)PLZ:7d@^I#39A^(Z\8a_EO6O=Hfb=/T_^<TBH.DD41BA[^A
MJ.31,1f#N0Bc/G2X1YaM=1L,?AXG^>UL>JC#c@BdVeLf.TBC5C7:^/\=IW]NBB5
2/NBceL/PBDU[efQG[EMKaS:L7faNP<W<5CKE8EMcF=0/RG1.MG1E/]8+S0<1bJb
ELSF@KKLBZXN;O<Mc+:5P]C\;DeO;?SFE^/X8&fYP(13ZcCMQI>^PdDC4#?XASd9
bO,fV03YfZWY[B^1Aee-@Z1R^R1[Sd6]BR4?fV&gLc6;e9#IM/LRTG8LV82=_4?.
W?D#Z5Q5P/BK)SN8O=2@5]\E>F/]<;1eYH)-M>#]82&+aOG/J:EGM-^TPf11XZ>2
?3-9FAYgB=4AAY44WG:_=_X08[eb5=<=-DFU)EIQ^]CB95JKTBJI0R[g?2>F;F)b
9&:+G_Le2ET+>ScD1;?3YGVN<6.L3D18e;W9_dF836A8H-;7AJGR&;K6=bZM\CSD
d2[9#WJ:BRQ1P7;a+)PNMID4^C]RIT0aA,7EU1ZW+YGQSO/(\B;).U1YY;AXK5Vg
g/Z&;U54T1J_0Keg)WX0]U^<6.@AgS428NL+/H[+<7e@E4I/2^dEbVX.XeMC2.JT
L@,ZVEa-A5&+[3,V6C:bBc>YM5_:1aXc5BQKKfTM&8&UKeY50HKccP)181R5AKc?
^GcC\3Vc21R8BZCPR3_HSVBYT07_0CG<gb9/cP:7fA3_MN@Rb(72S8Y<M;IAg,#V
b[=T@2GbAOLH06e-,adH)d98OF#9;(fM-L2UAbZS23c3+^1P1>HKZ:#OKZ].+NO:
d+R=SBAc^eSG+ZaA<IW8?\&)N4N94d7?I2,db8,JKQH9OUB_E5G:[eXIdS39+TU^
LY,/I[84UH4ZPcG&:H>;OY^_+W^QKR.H@ec&DK?8\/P#bA^b>bgd2KF/2D=e@<;I
.K@R#:PYgB_\G1QTQFSK#TXK<R4?YC&?(M;G2=F7Y\M=F?+]QW>AX]O/46FYZ\BR
gNK)Q2CcDSJB68NK,C_NFOT5@ae:_5FH12;K\W2d1=-]&NWZ\I-9WRBa7deKaeg1
Be>R1Q.4BT,QG#\e^70+FZ?Z+5ge,_0a:BFc\5&Q:&f0YM&XgbA@XC8ZE6f:#?HP
@TP[eK?H/QL3A)MgXaT(bY)gSMK@7[59:\177NB[-KSTKWZaA?^]dCJ)Rf77dSUD
=5(a/R^g81O)3/[L>R9RgEW?NB-G^OCaRaOe/VKf3IT+6+gI).Q(QPb?5_\H=]QX
EeKD<28:dRO\Oc]F7U)/2eP2<_#&ef4(Z1>a.H@,^3V&aKHYeFFHg?dF7GV5_CZN
8),=R3Z+9A)S=E.FgI^gX#cN;.+&KcRgO5D^R/]IeP3Z1R?8/HE/KZbL0\H6NYR[
_VH?0C?XTBH[70GGY+KC[ARa_2491gWFIB/:DQ+SfKaWS@,;=YE\+?G7a\YVMB-#
?##D+0CZc[0JHNWHCM37:1P;,G/PS\4#LP9IC2LLa3\P5c5SgfN34)&>7)PKB]GC
MAIRCdC(__ZK_e9A;Q3?44GR2ebJ8L2A2c-Og?=<NDJ3GW^<RX_Xc3MJ?X[WXT:&
8+T:2JSU<QGI.6NeENFDWSW?aE:Q?S,b2Z_7[gAEE;fJ_e=#.;ZT3MgO]e#fAF(c
RH3O>FE0QO<;G#I876FFN5SH9g-APEcQX;e-FK:E,G,^SQ1,:S/aX]BPaB8cF?OE
_IA+M3HQ,1<3&eGX+20LfBMaf)#943HH9gY0K04bNHLZQ5+=+5).+Z1Nb.V,B<gI
6(/G7@E#NWC[5<36cef6(U6W)];W4Z:=FYZ&AcHT.>.VAI>Mcg5P-TL2]M#QTdRW
^B7H]edOb0R?>[R-6A?_I4g9FeIAS<VceGOHHb_)_5)-F4O4CA9Y,0S\F1@\QUUa
98>87gT_TY<7NP&:-_3dEQ]#ZB5Ld0J=&AU3cE8+J:^Og8&Ie&3MSQ]EVJ5?_K0D
61;XHbE:L3.>)Xd?L:#H#8ND8.)Z+.AYIF>NYP@IY[\BIe0ScF)3&cYeb,8J;c&N
DEA6B5=9[8)@U<L2?db3:c0dNH0M&.c8H5&KGI?V]<)5,<RDeA^eVLbLFF5O2ZQd
4R?>9;)(,2#0TE37OK+W>dgQf_1O\)0.M.TaW<MLM^B,a,5g_(D4Z7^B#b-[Z-]&
TWTfeGb-40BQ?UE57EP>]<O^g@1[V5&+fO^JM]HK4N-c@,E9#>4,J-2V]O_<AYNJ
7YCK?2+#A)IPV3]:D]M8=-GU:BIRGHWZOD+&geS=L)W^ZMJ(BaU:KE[5IC6\X/S9
XEaK[E[GK12[>8IR^@JQ:R+Z,K+09cU7BKV>\-E1a.FeZ1(.T>9>^.0S@P9EJO)e
NP,1A.OKJ<]HD#J)8RXWMLIW3BS,c<3cF-=D==VdX6H5A58Y/[WJ@@THLZDH<@0O
N5(:OUb&GGWJ[5g]/MR8d^SI1<\ZaY>dWd<A.\(ZcUTNKU]7::fW##GCD(X0aQ8_
N2aG&HT=egCUZPCDPfa\6eC0QL7D5g&#]-N._@D,WT1EBI36?5;8IFb.-9,6g5Q1
[KZQC3]Qb6YJQ/6M;B]BPNZ?04(=NAL8W34IF[F#d#QLg\/be>M;-,(MBd5H<_5Y
@]8,T36&c?STN0TB>JC=7D/O5^]BK[3@TZMG)U=L(4bGU32FVgac+HLB,B=I<_0:
91Od5g>:=X?]N7f+c8+[RdQd)-(e?<-e4).&O^-SXcW@TFf(MaJeC&c6VP8.[7FK
^TM&_0;JK1KYd(/A>;IO&WfI2#M]C2<C^]L<Y<&)K-F;Z5?aZE+2/Q4=,,SN_8HY
Q6ac;4TRYKIB3KN[+8O_+1P/A@^6MM9+95.eG-:Q@;/gA_#bKf<U.G=(K+a6IM&a
3>0,,(.\SUZLca?UgD8)F&+g;M55=c.)MeM3U,(H\;;@K28b1d,^V)^[XOe&W5/R
[ONaD02A/P&)C\\V5(S32,4L#XKLX=WBb]3&1ea]f6MCV8>YKeH?V8VMF9Y^]T+_
&^>2&X69e^:B)VV<@1OTDW1XGb5Af?TaeU?>M+c#ISSXV-TFP=+P_6UagG,XRC?;
NaNJ9<a8&8fKNX#Pefc:fR;0?,MVNI(K8[B0S1,F]Tb;ER0[6VQg-XN34(gfKbHg
(B4X,ZQ<4gagddW5e;FC9:IPABGYQ8N9HP_E]1?#:?_A>JCF-DVL?beV&/+(86JA
R2DDN9Z7CUTRWg(Fd>6G/0@52XAL@HADI1J7;H4-f#S8QYOc]#LPNZR2NfGP55TW
6=O2>6b.GJ8DafUODC/gPF#7,J<2C4V[>eY[DCb_QJU4^H.BCVK0Zb]#+Z]4K,\B
3)S9237?]-+(_PQUTO2)3B\\4(8&<^aa=ZD/F,+LGe_I99DOT@cIUECf?02KXVb0
ZE&Ye3YYPL09R(0<f9BTI[JSM>d3PKY9F2#<RYcg+HW=IPYHB.6YTFR]1b^G(PP^
JaK@46<?E?QW\;2;T09WE02H<\_3MK[XPF.MQ[+Tc1?1^IHKaaMCd,9+\dO0cRU/
N[#S>e_9c;B]O=PSJ_.eCg+<TH&:KV;ca6J\BC+[1Y\5/EH3>QO3+C<<AEbS6RGE
=9Ge^IQSLRYRG?,<OQI(PeE@^V2:K?A.)]GG+1#::1NYV;VF5g_/EZ\g8UXb(,[#
R/@_P=c3/73/1KV@S6]T:YH6SIW2&VIbY7ZU>5#(2LgEM=-1)\37I.PHBg:6f;GB
H)H:g:Y/:#.;Y6e<B,cCT&8UXAF8G[6Gda6^K?0C8DY91VCGDG\_,M;1]P=fFW@.
:&-7XAJEZO#CRCCP,;_)Fc>QF<NRb+(5W#?UKF=JO9T(YNE=0GKZd:T7PH3Z#PR4
=O;O]6_H+M[,-NL\HdO>(@?)b8KR<gW,NTF0S&_X6]O&@c^7HZA6OS0[cXZ(IJF9
YIgSIPHb+88[]<YYW=cc^e\.?0GJ3V\/X7_)dd]7CIMUG&36K?S=27FFJ6:HJQS)
CgOg8]N2B-C[FgVd6,D#U7<5MU;4Y2B(=UT3::;L/V:AbJ2N8.c45g;JEK;.VSI9
X:Wb&SBTb9)P2U[^fd\\I(^=Tc#a=#6&G6LC1:D1],GZ>)7MX]>KTZdL/<Vf:(>F
7YJ-Df/YU@:McGO[M[46W_E[XA9e8ENA6YD>9P&(H1b(L<DG^=a8HJ6>g0JYU7:<
-PG=fFIQ5W.5O3Q-P#20O3g]7GXRed/8HDTGI6f488CX>dGKOQ,+@[&0BJ/I2_)U
b-A241(ecQC2?GdgJQM#dZWB&PE2?.3^a^;I=abML=UYBSI28SU99^V(=\(aIN:<
<N::g)Ebg66TV6/4eQ6]KH-Ha]FQW@JAU#E30\^04R>4eYD4F6:KUP>4F#YAd0WV
d_aRIcP11;\OgN1<1(S\AD<:Db.)XN9I@O1-g-<OF-aB>ER8F,Pg3BWCg.N(Vc].
3&--abG@8Q=^#9b5PG::ZO-e9E(3[6]<H6#00RMJ=3C2S,U?RKK_#6HX\]IV9e6<
C7TIIA+S6VA;5L58-85XPDaW/PG;2GJMDH_V4CX-+T-;>dBd,g4B7O,Dg>bDO,c<
Oc#5cJ=^/eSF2\;c^,gW/=U;\4b(O]DG:U;?AUfM^[3)RAGdD5&L&#+5\UOf39Te
VN.&^N3H3D;M,ZY8OdC-3Pb^3^bT:F>KY]_:[?GK1:BSREGZG_[D.fe7KMXX-a+6
g\.<X(M9D8J?<R,]36+\e#ZJ7QE+L;5P@;:KH:?U+QNf,.RNf(:5U99\WW=KZPZ_
^/?@7aK/WZ?<ScbDBd[Jb:gJ#8_1Tf7e@:;7AYAIcX40:5[4f0/Ob+;TgU[=Q-NM
^\bLO.1QF2\L84X;a,HJE(Y]<&BgcYO&#TLMF)S+))A/M?B=-V7\L4)W4L&)WKN2
dR#7f_ET&&]05@eZUg_=^]Y-CU8T,0+?5bDK@83QK_4C,/2dCg>eFN)2]HI;B5B,
GK9e\6b8QT62O7N=?/ZKNK5?BGB//Iegd.Db=/d:F7b?9f1>A:)BTD,+N[Td-1IM
aIcXD4NM+;#;&2Ja:N9?YQ]SFYgV4:U,cW@C>;W#7T7HH41.Mb6A>X]0UC<ePBRL
;DPg(\^_c&7SL;g4(NA1U2;NI&98KML[L[]M[L\DdC+e@=V6c]@;Y3366.cB_I0K
EP?#Rf7KHEcZ:(:g:2W2N/GOY_cU+=X(I]5(O#Re9P\@daB\HUY<1J<9(?+W6]C(
]+-9]HYJ+[IJO@3Q-6ECC_f.\AL>@gI]E3+Yb8Q(e&6Md42Y8R0VAEZHJ?YH_ZO&
]N+)29<QG&&1_+@X+eXIc5#>9PI<KHQ#XELZSBgIXY8M?E/@aU#^1:[R#aU0Ig&,
QN3KXZ3;e49+I_SIVO?A8X?+^,H)7]9@+8Q1Z/_IW4J9.D7FfcS6eIg.M==/8L.,
0-f8AAT][,-6@V6B405A._fbJE^O?PW[&OQa@9:;]L/5>_e&)2&bAb2UKM#;8XN^
L^-X2YTYC2<@HaaM\68(?9K[N6ABR)R@Bc;X]L+-A9XO.567(gB0fR_:/@3cIOH8
)V/Q-FK+_K5-4Jgf=[)8&-beBP^Z2>)>M;Q]:A,^a6_+3+91&4cE]C.QQa6&a1<P
d)KgAN+^Y3=9+^4EZHPCA24_cD(31KUUIf9fZ55cYZ+M,c)V&MH+R^9ZL-)B[QN)
9E;(9(I)N3GBZ]W:G858>E-+Q,,YENNIYE>VfX=.D:R<FCF\f7f/MaX=HQQ\Q07?
1#0&><[R?2>P.)J+SN[_R_-\W&O^HI&K-TD3[O83H0K6[f2=dPY(U#&NWSbFE:K)
WD/Qb2SfGEM__0M3D4f+^4(917e&5VJ3Hff=LM,Y1TYMWJZ(NT3S<N)S/X>BY#CF
-Yb(,,+9ZLHVPc9[gZ[^D[/I1P#LYC1:LM+V9&<c;P#55?GEKU4Q;,<MX+4\E.R+
]OP/Cf)(HNe2>^X\PbN@f,WA[PK+9/BfF;84KN_5U9TYB>ZO>6:E0OVI3AHff1;&
;<eSgR8[=.V6B[f5RMRaSFZbZ^#)R&:H#a[//G)WGXY007QARNgF94.0KCE3?[=&
<<cB=?W._bPDeff)M;;8;)Jb+7L=6-MKVAQB4?()+e&VFdK&6FP1L<);WHJ^<T^3
W^5VN[;MX0e>I&(\0KN_ZM-E;;ZfT[C&EE045V+B5@4^1\_1MLXNUH50S4\2AQ?8
AZ2UO1gT<cbQ-[12^b0c6TUMBH6ALXVQNM=;QEM>^KbU5gB=GDS:YM+NHA?a?b/e
/=P?;bH#_<UOR-9T4(RE\X,35+[?;M[2[Mf&8@fT8TG-A,Z\^P>]/Te3POF>-ge9
]\8V1AM.;7;9]eaRC9K<(41P+9ZI4,43PE/-gV>3(2DU1?6B21cdTffVb&5#\[(Y
QM:P=fY9Mc<P29N3D-Pc?J\K3_\1KN]4=0@M@4^L]bBPA:aR_6Z/>]e;Oc10f_K?
eUe0B,e#:EUeQTE^Fa^g:YdBT/DP#M;RLbMZ;[M9IIe@=\BBaX&8?ONNM+=a_E<g
XY;[#;28\_G3N)#/:WQ#QbKTcU/8Y6:U.05H]Pa^<JBA[71K4ca^)9=8]gc1V?Se
Idd/K68\1f<^GDc+1BI\DVeQI<]dDDD2[K;]R2BM=C<[^AGOQGM-PU-N^?F;X[:D
VLQ.UV5-)Y-+ZGR3cR4Uc]T+;7:#D.)d.9#\(7YP,8.]V0G0^PC@eD&IQ6)IDT;P
O_B]6(_ZV/OI?<\AY.DWDTLH.bfgLT@0X;g7<2c8G=.+D8eP2fP@7SEd2f3<>0g(
0)e3#K3UdHFVY1^.+;6M]AL2<9V(<>B(+S>gLZ@G;-TYSP?#[^2d.EdaICA,eYEf
eLR=Ia95U=@GMZZ)6@?]6cECfMFPZ-Ge:1Ec79UfcJ,E9OUG2c._SMEcDGVEN5(#
]V5F?&<9Q?A4,@VGS=N[&PIW_]>e9MXHLDHBeH1WYe.B.b<9I;EG_Qe-Xac-I82D
gYC<9-2LHZVPeJ,3a^R^MC]#^;6WdI=?c82AaaUB/==b;IbMK\;MNBV:,H0<;&)M
Ic[R^L@FLd=b>bIZ1+-=C)cTYN03HS#&K3:YSV.@#2ZHR[c18]cTVI26/&J&YPU>
.gS._0>L2I+XA5-I#OUL/-]:/e2C#N[M^R=68\Z\+1FN46BE.F2MS)]@,^5SD#WQ
aO_5Wd6/e^g;KY5Y<=UX(ABd#P)LKE/PH&<4]BA-K;(=?_,>EQ#H5;8DS@B_:U\3
S?UAcA>A\:[1X_-R75E93S&(fdJ2)6P.LMOO-]C&e6O6.D&7Eb/]9WFWcd]E#]TP
\@DZ^K[_NZF@aT0eHLQ77(UF]0+_FXB7.(P0-F6>CQd-c2IPLGI1TZ+@Vg88W?XO
5V@5=JZ43Z,f2A0_4JR5T&FORS(2L>5a3:T7K@-1R)TcP>0E+E9VA./:-YYbcPK_
F.0MBg5d0K@Y)@VU&Ta>;ZRR3[AI]d/b[NRIMJ@S7Q-G]E#N0ZM?P.NLJ8Pa0b/.
M.)K8AT#L>QZ)W\CAA)_3e;+A119Xa6Y=POFN5/d#<EDg0b\]df3Z<TL;=>V@c&0
Q0,[3(<g1U\A(RNTY4&^O-C/BVagIABNQZX)/G<]IN9=A6e->RF##S@^XS7+]ELT
0P^5XFXgZ],_CYEVP6c/1P5d\:6&N.d=?=NUV>:^Mdd18C2bX#;FC(84LB#+.O<g
@;>/32)HX@D&6K^SYb_771a<BNb1XOE<:?J6/+#UCDWNbY#.7OSa4F_AAAUSTPM?
L[D6K&)MGcA6fOR_UON@(JQg[&P&\^WVKV)M:4=SY>DGG7+TCH=+PZSGb\J3SVa0
HHOAC>A\QaG#d/@:eYDB4,QF\6LGK,PMWJLPaU83K:2g^aGF.&-NI4;ObJ84b+N4
6LU1da0S8a9H497,P+Eg>5SRY1?4BP0PM#P3WK_6</+7S6O(eM82PF1e-\P+],2=
/T1B]9bW];B)Jg3N]VF,CU^\Y_GX4.NL;69^RAA;Bd5gaP+II-g@S^YK)-c3([O?
MM0>bffSA)aJJQ>/@H0Pf6.\DN-TDFGBMcF:O>5,3b]Wg4B3;D<#@)3c=_;E9O8a
dLV2;g8WaeJWWF9dCEK&3)^YC^/.H.5EX=S_M,EGc-REO[A^:Pc&f2>f0:>C7#L^
+cOL>0_9f.(P+EEGUcY#.6JXM1Wb@Y&EdO>HQTfcUGeP;JWBCOK6G?_LdMB(Q+^0
g/[EWNH9dJA;Hc^371b&,\__-DKE7Pd)F5O&>c6bNbJQ:QZ6b-dcH\Q^=e47+X1Q
H;f)&;#fSNNaYE8EQ6-<S^JTU(1622_4<\&.]R-ES5]aO]T4C[b+IDgLNPT74-8?
UU9dJA=&gOeOW9.WE28RLEOIIYZ/C2LU)ALLd6K.6<XRf\LH[2]XI=#P&M<RCG+K
/Q[[<51?F?LIC[Ba^aZ[U,_O,;_BF/f[@CHPG?YLL8U=O-Cc+34R&FMA:@FYU7.<
W^A.BfASPQ#3+W63L7JT>Y<I/ZEC8)YPH4?WMS)f,O,VO_^@I\K#)IGOPf2DRd]W
I:eY]LCQ3X(,J)NAgYTDS&GaV(R@59T3J/a;EfX)\KHU[]+R@4H#+LJ\T7e9YCH/
fRbG1=IA_1\O9W.FeJN/TE4P,65T6]-Z_\;/3c88G./>b(WYeH)&T1bXHCW(:JP;
\=2?<P9J7aA3;<:55\8ZFIBg<DHU4VB:aB#AQC)HZY,U.O]FeH1:Y;Wd\,J]YYMc
cLU?(gG0-W/=HN#ac@S[LeGcEY4JZEK3B>J^S(?cDB9fJb:.T.;?F.^K94-4=_##
ZAMH[+Q54c5U;N+Ae\G3\/A\K225/32-.T4EV66N_IRbR@&Y](/Fd?LK-dO3K.Mf
XGbMO<..6RJa&dMB95379TS?>G(6,W.<WY05O_?e[@8MKO]G1c=W51aFd25,[C9^
5VX1^WCVIU?J;37]NI,RDA[W#KgQ^\>KMRc6Ge;G\#8-e1-f4Ec<6/b\T(7;M^F=
W[bGZc.M<XJc\c/Rg1FY7ZaD@TW>K&:UWM#gc^QH73<BB;HV=8K37PUR->a5C3GR
bF&R6<MG=U-Rf8d>OBAYd>a1>Q5G[J>GY8C)C]TPT_N6;I]MDR0GafDD;H/H\D/(
A-J/Z5O<&@:R>.6fd_7QRZG/OgCFPb).BG?6I]D\A[IAGP+&M_E&c+D(NSb/f^D1
6ce.7BTT+PR1b&YF=K2K\&Yb\AfO:(&e;07)+Mb)>93.23+.5IWf\7(A7?T?A\J+
,ddD2c=;6E9WJcWW(:)AR=BY<)8APN8Y\CRBdK:ZE#B1J/aMDW@]G#:2bGD3AJ@O
M=+S_G_cP8cV;W&VF4@8B-MVP702WPV7HfI.+:,3HY_S?cH#H^_FOaEH#0E+\E\e
B[g8^KMccQ6U779J,_Qe+cVYQ.99&>&SJJ-QG@ZR_T]QX9,HC/CXG@)Y20;>T5J7
\KI6#Rf&+IHe?@O(P[L&ULB7-Wg?#fWK994RZ]MO:^T)]QN)7?aS320,9Y#DXDVP
0R3eQ5JQ(dNS4a@)6HL,gERFcKW#UTZ+X96</FLcL:b:JGMAKC_?V(W9GcTO@B<,
4&,-.Jb1ZK571LO]g)B+X]GKK]5,.D-&].dU=+gQRF?ISI/24[Qf]E?5fI;8#+C#
g_TeT:D&2XSPb_\[)XL0>R;Qd/J/I>/H]QAX_[^/BA,J0?OX^ff2>c&T0dG^H&^G
\4>B3:?HU;)cWeVfG9H,:ZcLMTA=(^)+AS.F-@^;@>ZA@f9M;N5;_SBgO/?=XA_G
_WV3dQ1<WFYLZFNALVf?R81d<-C6:NeJA<\d^RM+:SOAE=-2+2?Pf8ebJ&G9cMT=
(<^b913^?WfB?;FQ21Y+TVfc-5/dVAd73C.67;[][NeHBZ](aA7f3VQVbTLLfM0+
d;F7RKf137RSK][:-fHG^2G??1_/2JgK,JA4?W9>2L22QYVK],=HUO_SV#TK+9.I
9DXfV=AM,&O=D_(N5J2=aG(8d5VG+a;.(Z3O8=RF>9BS>EZW=TU#JM,4LO,gc>7D
O>D-:cbQ,.E\+-f=&WD4ggdPgb@ZG]Ud/1HZcK\K29E@cSV@9X3C?14.-I4#J#Y5
_CRTF#CX]&W#XO4T-0KQD0->GN7?=RP9^>)c87]SC<BK+71^eZMT?@6dPg.Q]>V0
B\SRV+4F)PA1ZJ7NGE2aQB77WJ;?UXY<R&Nc#=>Y?D(;V0_aKcbQ.Z;FA;B;_&;g
MDU]IN&3G^a=L,8,)D=7C<CMZ1R?S:=1K2>Od8[XYEVBV;4K-O08WYY9<T+/c0f8
(UU(R;&3E=T;N5+P4)\M6K&a2A_,aJ1@T[O20OT399H+K0Y/,Z(ZaHd-_4OSAOT4
VENGe-A-/-bUI<=g^L7GS(\@43S>e6]=;AEU,G&\b[d&?V)+I[TfP-TPA<:<eC\B
3-#(>&@@FOd(&b=?9Yb.R6##BN@J&,\2LHFRd>=:MW7cITD>8@@;L/7DUS3^DQe/
dC)eG]7J@6OdMd)>.L:)J2_+?_O\1>;5=Ua^=WcZD=]4<E\\H7CZ(f7?c&7\@^7^
EYH:3#b1CMe=L\D=RQV#6Q1a+7g-b[\/5E39a3V_P&Bf5O?:fc5))GIGK:SZ&JD)
+T_Q#,<T_c[SMM:^1A/@PCV>S0PK(LF,<M_LAQ?(&9]ZY<#DTD7N;<U5418e1C.B
6Q?@[.f/H+cUDDOF]#ZHP-dH>M^Z@.c629Q2Vg#.ST(I2MX-c3.&UcOH[GfgRIDS
],8XT9dGCA,S]PE39fb+(.fB+:bGJI4V22,00=HeeI6SH#:.S_SLU4_RJ40A05]@
?UU0&-\.E4>&=8DcY?bA6^gg6V.U1#;PS5d(J]_-H.H)]7K:H77YD^=36;J-3:[7
GD;=</-(ZK^85?9[2dggZKGD<:aZ)9f,gELd4Qf,g-Vg>KL]3LS9=,X/^-(U6eW#
QH6@23Wb#Q[Y?>dY@OXFeJL1Z,Yb6&OTd6dS8_XA6F3GE#^beQ1\IR1R_17L,C]d
:[b7B,]9&CUfHQ5\FV6D9&O1Xa=d]16C32:D?4,:XXD7L;R8M_f?;X3O+<[YaGS]
D:I7;\(g8@^Q?N.bYdQW=UgJWXd#8VZGHTLI3DCCDQ4_2W7V;4F_RG,6#]=S#(e#
#\Ke3?AHd6^b]H;.L-@A(?._NZRcBDRGK<a@8[dKJHb97Q/FNQ=[bIe\=DDM_.W(
e,27_-AXLd69G0P[\ZD?1SJ>32Of\;&b-U1_EEH@eTA\K1#Y+J+cQLeCcJ/eDDRE
CE4G:?B,-)V582)7B03+Y>9CY,R8dg&[0NFWR(HH=gVV+T1bfT7^G,#M/6D5@JcL
S,SGL(T,8EgDZZ-3LC^0+A>3Xf(K,<Q.2\(-126=fM=LgEFbP=7bRG@g.I+Dg9T:
f8S7<Qca4d;\T)ZRMSC(5&=?U=c8D5-b8._E[W4.S(>KB-\Y<LMEDcH=2^&HX+C4
)/#ZVJ,HZYIWWL1_(_>T5AY4;EH:82>?dK?LZ1eQ7GHJW95+?HS0#UfdKFEI)08#
K88a+T^JIO[6+^7Q@8d[[BTP&U[66ZN9,+ORWJA?Fg64_8Lb76PXK3Y+MN0#/dE4
WDK,[2#J:1]T?Y]+&ZZ_1CCe]AF/R8Ig?PP7IL^A2:_8E^c?_PT_G+Uf=2G\?ZY:
HYS0__/3>J0))98TB2\OY3-CTJZ1K:4_W5WA9:C:UFA=/RX_>;@\]00G2N\dg.fY
bZOf#7Y&E-(?5I/CFS&)LQ\J]#+e-P.^:S8d?K/OW?.A@I\,IGZ<><P-5H\9O3JU
aD1b66Na]-U_e?&eP.:8bO[_EKP#<TPGF+F+?>/B+HYG6S1P^+<]c+J;&@MVV;bX
97WW;P#\ZS9;F:A)d.QKZF#YCJ[(XDg6AV,=A[86T:.C+G:V(D&5&<DF+.2NcE7g
aPRNSQTE\CP5:-aFCL/-5Gd4a^T37I[L7.50b(MfJ53_)+C\MDG:>O6?b2M@EEdE
>0P-=HK1T204?3[3@-gX(,UYaJ>UZ1H#a.e0D:>24IN9fZS81)HNHTIC1_FcFY@O
Q20?[SfI8?X:eX9eU05-4SIBLF;Z,GU92ZC9.L?^(bF,TF;4A^3,>YHZ6TJeBY&P
1>#]?RV0]bGHCQ^eM?Y3DEL:AYDQdM/e[?]&#/T8IF#W?eO3)GWHEb-A0eJ>=@@L
4BP8+2A4-NJ<B#[M260<[&2A6J#FSgVU?BIXF158fG^U-26DO?HAB,U/cLI[SQ-Z
PR-TJ)d[WBS+.B>-LSG9)T^YPF;aQf/V]E[+M)DX_6G4]7C<8;X@-6O9Gb>D=[+-
GVOcBW;..0>(50Be\b)ZHDS#D>4?0JNRZE7Ke&AX@+c^PX,Z;97d/6Z+@/&g(8MX
fLAC3QMSMb,QE,<c5\O\ML4a[20;JVCT[H2CTSc;IL>D_E3,JTZA[7c=R[bSNAXf
N+gUB]SCAGAG;=:>3+]6cWaPdUIPcMgO+NG-7N_JT^5ODL2]YM=[C.>Ia:@VKR^c
+Rg^L2=:fY:P(>b@g:IgL&Ea>VI./d4>)aJcc?L@@BHT^GZ)aMG3N&7NH4:P#=3e
\-&]M@R2:STD(fP2.SEW6D,UTMBNY\X]=g031Bae(ZN2Ad)[^G?SJXbE)d6QdI9d
5.Sa.YU<1]:2:@UOX(T#92?gK0T0CN-7VER@\U2,cM7dANX^Cg<;=NP[.9W_NL67
18e2OfcCb@E#78L/E0;fN:ed:OeQA=/=H_#,M9.;XF7KQ_^K(L8JI8FLELb/CORH
ACY9ca,aEXc\7gEKSa4,MD/1#WYSHE.L:X?DP8=dAZ0]-\F(G<95+c9f00@;.35>
V2T&ITS[=S5BD:9Ie4a6UKCYX#[TU<)5Q9F>@,0_-O<<0)dV?BbY2TM6eE>-NX7P
Nf1XaB8E@353aW328NQRPV;aPY<^#)K3S,gKM3D]dJbBK2WT#)/)S_^\c#9@cCSP
EZT_&-4a7?OfeFXd[[1O(D3O=;/M4QH+P\.A/O_[GVD(WFB4K70CS2GaBc6XBZCP
;FY/\^M.#>=:-F]0\-[OCAVOZ-D>T^,KgF193cQO(>9)J2#CKM[NK1B_=6>6T.-F
(HGCR?g@fM9;/c&.VHf88?#GV,O<N+M1]._EgTSQXOB/f.GA#SPbCg5,<,AHYaC&
Qc:?RBI(>^Z@&\B>B9QQ+a/9NQ27]ggUUe:g(8+8M<3Mb1b&f<XSM4+?S^O40(F4
69V)U1]Sfc[7=fGBbBSWUN)GDHPHOgJOTU@_cFLH8O8@M1VC<F</H8fGJE8P+DCf
C\=CL.)^3A<Uc:c.(>8S^)>W_ggYf(Ug=\cR\\Z4(FHP\<JF&.,[CZQ.I0f39b.J
PG:7#S?A<QH@V=@@+HeQdN/8RR;P\HAQa,(bY]L>&fc:U_U-^?C&e\F2<5GW.9aR
L<U/A)LYEcT51B?DO5ZfcaP.O9N;Y8d>adXRWUO(&Y@(5=S]>L\(SdPKRbaCS(2/
1Y]^3&WP-D#6VQP)9beCW>#^>0KAg&Q1;:B4@B?:X/Sd;)]dP(BUCY1dGYcdUFg;
=]GR,:gDLK_?/EPJfMa((K+MV<JeIDV=X?LX(ZVd12M/NBFD1]1=b_,>6a1YP(]A
]B,.#@2>5\V]AEd_R<<RbDCB7SZ/1>KV?EHUdBB+Pdg6_FNBSM/#(-f/HX^>P&R3
EOD(-2?)=8b=1;FAaTKEJOcVX=+@,+YfNe(g36Y,=X==8_4_P#V6Ve[//H1@ee,>
Ig5;DB43Z2a=Ua:V6Z?/LIP3_dIaV;J>KC24=SfNQVMRVO=O],+UO=8DS3U4aFAg
aUT2;6:6\H_6MKbI>5S_gNf]DN0#dCJ38>0L]&OCT>JJHH^U0R;^GH\QD@9F3\fZ
DeAMOGH6H:S\_+YgZD)Efe,>Q,d92QX17D121-:-AE@V2_&W2E08A59H=X+=Od>>
/9H/K8K/;A?.?KIdI5;=_.fTEW.+b04TF&,RX,29N-_Ua^0Zd-5L+60-dU?HgeY/
HYE7-JSD_L1Z(]O?1\7ZB05-7D5VF9&:dRKE15MM@2_UIIHA<1J;\c@]\;BXPFOW
9(79@8QAI25=,2bcaT>a:SW&)W+Z11\\<<bGc_=e(6IFEH,aK1DLU,^=(.9MYF1e
YcTac:?FA_AAH1ZDI7\\aQ7=])V<^fd4\N.KAB[1-]gA7?LLf9>d,,aP-[D/T,f6
bf[-Udbf\2gb24b.\QUcB<1bXHOFYg3V#7J8&NTd5<K[dA7#L)68],QZ&>(,[S9N
:L-a.16_35:^4YD<WRXF-V<^JUR?U^]fJ@JG+AG^]+4.NCeN9d^\DP?JG;aVVL<@
[@0I\-97Reb[Q14SXV4#ObH-[\,F.eLfTXCS]\7=(aKLL.52+:b7^OTNf#bd/C]J
O5UA6E_PLe@,W&&4]6M_>U)_30IU5.FM+Q&L)P?4,.[Sg_1#_\KbN-S>-g8-:F7R
KAgK,:50LO86e@R33;:@?4cT/V?2/&PZQ6g1aO3752:eTdUOLeaXF-A[Uc-^MfeH
:HS-OTebNfZMe=9J?&=1]YS<UJCRM=UL2FN8[I_8&a=6J&RWc_T[LF@LC<99XTCN
8Z]g35e@;e@NdS1dA)VHb#C?b)=<TBbOBMZ.^OH:7aVW#QM(-EES>QL@39>Ead>U
MID/1+GI.>CC5A<,#^geIf\R@cZJ&);_/;<;8Q.bT+dU)e#g(<[B=O]P3&JN(S:Y
.f(2?:UTVQE9MVg?Z23#.INf?O^eT-(?1M_R[Rf.:UK3.cRP3T]9eQ/YDNIESRI.
XfRQ=NH(A6;6d71(F_X#=[6/9)ZST2=UKV&6<>E+D=H)&UR@;T<WT&ERID6,ANNS
<[0N?12K2EbD5:\&g2dNUWg,(4-N.J>HWCG&eL5863FOR3P9CPI#O7TZ^W?H/K6.
0-NL/.f5S\X1-FY.Y@E]+G\9K&CVWG&JK3Z4&XPS^ZD-)6fdUZXJU5EAdf.J4_fI
X+YG?LPA-07<&Kc]3E<@J/L_[aD,<bO9e4NA&8;1IcA6GJ@AG=#\01aTPM[Q]31b
91B?Ud8IYR7JM/>^^fcG2M^cRC=R-R+)L)BDCZ0TVcfHX8-Ecff0/#9a/R+SEET\
;8VVI(BFCN)9(ATE?Ag8\\=AUIZa:/Cd_9ZM.KJ9P9/gBQ)BQ7KCNO\5.MFYLJC?
Y-NLbR;@D,[LP+N?DCBEX]Y=_P@TaYQV@+&OW\ER,C15DKD3?XWDLK=Ne,;D.K6&
8a0_.SYH=/&&P0g?T:P94U)[[9>+53N2MP4?2_7WFBK<31L^1<VMC;8c5M7X?[=5
d2V#B4P]dIQVO&5;HX;+8;[?gJQ<=bJfQH#]MKcJ?.Fa6?/2URLWVXBb?2L9b(L2
CX#5d_CXe\a@c8KC#(ZH0L_?g3G[5_S1cOT__>f?\WETg<A_A/5daNZ[W_A??=.0
]0Ye42Rd^]:.4)_(1_\8D&2geE.U[)RID&Lc(6I9B:g\F4X0^P63=5J[F2cFC>3f
A[9G).Dceed2=[KcbKSUAVVBB\Kb/)@OOeQSC46=;bOAAc8U:9KCgA?F.#cVb^M_
]TX,a]Tg@Y+VeI+Pd@aD[cMS&?_Ng?#NJ0+?]:f-,+SJ?TY1YKOc>9[@CI>Q[[Jd
D24F-AQHTKZC0A&#.,CL7bd-)WW,_B?V3d:FJ/8Gb.FR^9c8abKBBSRT7dH-?GI_
I-^L884K_5Y?A7E1GV=L\c<Z@DbK(N^TMe>>HQ\N,XXMXdT+Q(0g<S:_P81McCd#
R3HD6NV4.ZMgX=LagdTBK@-[/CYXI(fPH7aBUcS_ZfC<.QDe(>Gad-YDZ6,4H]+G
OD?_ZObNMVD6@;O)<@CVB_;@,#K52QG[^S7f+9V\UbCgb&<\6Cd5Te&bTA27^94D
G>c3+EM8,3+2egdWZ:3H?J?+W\+4(;+.\4+\fa9&3dfSfbW#&6e3AI?:^3E,cHBX
Q<PH^5UfINHCCVGJPDcdIM[?/Xda,OPcD[.XIVb]BW5_FecU?,O;\:HUAEE(c)JJ
DX\M,b)GBZcTZL/Z56<8&P;LDV^[.fROAd-6Y_&.R6QW@;c;V]J)1cUBRL.ODSd6
VN/D7B>)DQ2g_aK4_NXa[5:HJeE^&fDLTXKGI:,77/L53W]PVJ>3aH?4/9>NY2SN
X4J>e,1bH).CC<b^,3@[-dQ\9L,(eZW5/X-32TJ73][-6XXTB-G=GN&HVg3MZ&1?
g3^P\ITL4\a6_<d@ZA3ER;_.#g(7JdA0#bJ?,Vd@1<IH8VF(aU[OLTVA4UZJf-WO
:]<F&a[^];]E9DT4=)5A-.Q\Y[b4=dU;[AY/_.U@AV6H/\D0MF=>U^=CMAQ;eDSO
O8)aAEgfXbb7eP&KeWJ#H-YbTS;4CJ(T8<SP[>CYLXV9CH15US\#SJ3^N70>604Z
WBYCE:G0U_2Fc=_eRR=N8-NVb:0-3g<?.?-;GX?b-]NMfFB/C(8A#;=-a)K209B]
?O0Ifa7<KBMHe(+OA_a:X51/bd[(Ob(Q_4?-SW:1N&8gSAcD=Y2eFX]VX00YMPQ5
C_F>UU.a6.R[MU_=><+\aMM#1Ra#B?HOJ\CK?gcF?CeLK+bQ=[@-#O7O)H_G+QD?
FL(GdR_VHE]0O3334NZDY&FG74\MV20?4Kf0UI@?N?E<J>cMFKZ?T\)SOBD7?\&&
@[V7g.IUFZFVU>-0;.#/&=Ka[YH(7)/M6E5UOBQUT-6=M#@4Z&N;BN_,31_5MA[b
.Za9>=QU.E\YV6?Y4JCa/Fa4Yc,:0[<g1\SAAV)/dcI]C,gP>P^NY>3#\KgNHFN8
M>d@A94;5I3?(+g/FB:)WB3W;(YDcV8.[WfaWQ8\NgJ]4.?b.A801=>20^8/CI:4
H??+^0YQ\_RKA8eEO>3LffM0A\IS\;)I03RcUJ0H);^FEb>,>?aX?2&;V2WR9ae6
2/5\G#)&SD&<P;+=CQ;a,SVP4L.4fUgG)4HbYg9,-&:JJ@_7?97WegCT[Q@-NA7[
JHH8GI-A^&LBc\,D-a)LZ,#Sa9E\JELT@d])GR#[IQN(8c<K6=OF[I6dEfa?;J3R
H[NVf2aeS78P4S\XZV?;]NgA,6>=7QM-/B73e00#L-1C,LZ6::HeI2ICNLQ9Ob[2
+<9M8XP1M6?^YU\9ZVXU0^Y5,e0F;<bWB\?bD[S0^aRCWDOc4BA_KP_C-9LQ6V@-
?FKEeZ5\@&CdDX[#6&VdDF_Z5P8B/.SEPX79<eO,]W_PJRPSO2U4Ae-Pf-Z/b5d9
-]]^Yb.=42UWbOP0W.N\HcR[=c.ATJ+6FfBL,0G;f5_W=)91bKfF9\BS:Jf.1MQQ
D6)1UQ>-g4H>\V6T;)6BDOIMO/>fgBC9AUU\OUT.&6A+^=IR?e59,RFWXcGg+c//
I<aJVZ>C-X9Q8.2=#VJC&I]?;#^<]DY?Ka]]T>8&D:6?&We]7SWMGZ(e7>AI/S-)
^SP)WV9bHMB^U_JP3R1<W.V5^^__HDJ\XGRWPWBYF6dSJA]Fb=aK;YbG61\\RCRM
&#(XcB1N4/5>1R^>)>Ng,RPLLe_QUIS#RW@/)]a@E>3cDCPMOWLQF[USGAYDK3@]
<1[A>3;2:Q<aEK:80aZ3Td#XTAOc,Ja_^,eDa,C\EGJY[=^U#;GEc@[d:HQ:0@ZD
.T&V33+\W)G?<PVM+^6g/aG#OC96__L=4_AC&BJO84C&+<XIgcQ/N:X&TXJPT\2J
&:RU@O9V.1Dgbg?<W0+]e=/EQBZDZ+de1=f9J_&);A<2+M#\B-W8&[8I1R+)074Z
_],-H@<=;MfCC9>Z(JF4QRCYR>cRF[1a.;MJRMZU&75,JY[R,^0=F[RaZI-JTe50
GN-Y?@QVdZC7+S6H0d72]GNG.H@K0a,AI3c^]A7XM^V/HSE..Se27FT?+)A&]A_(
;dK)3TEdT&aK(YLf)P+7Q\31e@29#8aD8?8>L1]fG=4T(6_B2Ic&B[_d#Oa9^Ja4
f\21C[\_5HIVTPEG5-DYT#F3(1(H7#)=:<R=5G+aEAN6?Y-S/T036-K2=44=M7>Z
5gWXN8G=2fEcR3:/#1WTNBDcPQZ,9Z8d^(K57fbOdDS&1LU:)Uf4_#4IA5J^K\9c
>>[K>CPB>WIX>A@d6-YK/b0QQSe,M:Y-<OZ.9gF19M);TaOfFD>>AXMVSeUUKSJ<
Ne@TV@X[[J7SZ<c];4HZff>1.P@52.;-d8cAM##Vca5/9)M/RX)P=,T=GJa\II4P
+5D@>O?g]Rb<3TCP+&KB#/9_<HX?K9STY3MM#.0)+b3F^T<?#b9<T2AZ@WN<70;3
?>B+?B6/g6V0ae2#,I=W54[TG4;U0C;^Z7Kg\6C-QL#OeMHgee)C3A43WI<CR+8P
C)4UF9W-89/E=-C8a.^(U@]D<)>d)9^e3MHcP-?LN0LHSY+T\JLAc5GS&e9=5BO.
GcN5b&3JG#=3>>:<\eRPeI)H1((^X@)]#<UV&39:+156eF?[GQ#K.\fc9b<TbD9/
_JLQEP)U[gdCKgag3&.)S-Oe3#^W:-I/Z8XUOTT2-JYOK98+-6/+X_UD6>_X3:=J
ZP8(ZSSZ3Hc;S>SB73\&)Y3N4F2A)5#3Td\+;g=XZ+[VUb-+<M#SD[.I)0^5,VW3
>&FGb/,=TE+S:./\Q;;f-8#TGMUR)_]I[fZQFWDSQQGYGaCdK8>S8.XBZC-V7d-8
BU=PMJ59EH]cG8G0<:QIZA2MbS#?CGCAV-f\GB=K<LdHP:UHLg<KK3\)W/8I057H
MVFXfG:#+2#Xd89UT>B;<(b+XL3Kf,P:[cZVNZ+EbXfC^-[J7K&#->eYG3+RXG4P
JV.J33>A,]N^_GZ#LODEPK02Z.ISEI/MWUA=2,_R]]6CL0FIJg#?Z:T.27#T)X-0
QB2@?+0URU-6G^J[Je.>e]:VN^f^,)6<=4GN/53]XG<+K21eVZYbcJKa0NJ?/=C.
NWSW0Z3[g+=BP_Q=,V/?9-[L^gIL]RV68#7ZWeGGPc3R[(Oda&a/1gEQH55cTN].
I8e4-/Q(@Nd;(Y.J@d>]a8M8M+-a,b_T)Q8f0;KTH<a&#g/O^JDIY>XFX;2<G982
DgIWS7?J[.3WAPO&23HH,P<dX=,I4dA\T0e3HPM<bKfKFSU0a8#AGcaOR0A?0]SO
UeD<+4?(ZH:==C5^-Dg#1T<&FbM=ZD^HKc^O?N3S6LN7L:1R2VTe>^Z[/<&g&4/Y
PCCY:f=c?I;gc=R^Zf[DDQKXE0dAFMMd=LS#=f4B3fT9UX>@-:SNEc#,OLP;Z_KA
?f\QPCceQ)aX2\5NaSH()HHFN#<\/Q8f[?\[8F6I(TI]cE7QY4G\QQ&J\D.YeES1
R#EbBgP/DCORLMTKWA4LM(70O1(ESO=#F5><NPM)+TD6PA2+/5gC8)LB)MB.-:)E
6E,:HQ1KdCHJFC:[;Z+cOTG[-RK>cPa)e3V9<CG+V_IYG:KHUIYYCGOB_NHO)[/+
B_7@TXBR&Y3e:XJ_a+#(Qcg?=A0\Ne<NHE+F\J[3]\SXOI^F1f;,35:B3TN?EI(6
A.[#4fVNB2Q&&4E(0BfW,IUTVe#A]5_gO=.c7f6NLS>XJ(Re9K^;MP^cY)4BFX;-
gC,6J1dZY_?d[5CAe@,dLM1\=X=H7?0S8RF9_H&[;OH#_\E61I288<63H+K-[YZ7
g+W3bc,bVb\+2(8Q-N(OV7P?N5BTXQaYV4bd@6#B#O\8M,JWUBI?MQgIeGTSA8g3
XN<XW8ZF+ZO\GKP@)U(VRbDS2OF1cK(R95?5S/ab?4eOQT.bTU#Y[(K>80<RY\(Z
9R6\(bVH?DLTX-:,-@L01W(5:4UPUE)1FIBI1N/2R1SO,6:V6]a#.e<L@=T5ObaG
)\.,H7#PJ-]A09626ff>)^J<E^?;9g0ec2&IJNN:NQeP\I1?BBBXF-)Y+WLd0#+5
EOB.e+?eAIS?(>YA@.8>2@CB]V.VMU#VW_&a,[,9U^XDK\<XaC))XLWb&Rce6U<Q
H9?&#HNDYS#(G-D=5A+NS;2+G60;M[=C?W@Z;aX5U(,HN-CJWC_&G^..9?Y)H1e-
VEX;3[^g6CNHA39(F9?8@cC^[;7\0^(O#/Ja4@WSTg#E4Md^BH#0PPPd6=9c&DU3
9ZePC25]7O_-LJ\4H4N@CL.P0LB&MZUgWL+B)B1\\1IIbdc-:OL\2KX5Z5,VEESN
M@=-0/H(07=e):&V>VQU\IDI_:Nbg.NN14#S/gFY9RQNOX>;)OH[JFO6P(QY0]GF
-XY,=[3/)65=X#Qe.>IBV)@A_Sc>CTS5\+E<c6IJCBeY:^#88B<&2P[3X.fSDNMa
HF\K87@^)Q-#JcZ;b<80.?:gV+LRb^RF7I4=Qg+H/>dT0OGB?197=OM-4=IWPZ#V
F8E8;KE27/?GU[><MLH?G_ZLeH9Z=a(73S[(-KH?LEONH@O6SIJQaJQgFJ\ReBDV
^RdG<&fJI,C1OC4bQ1&X00)HA8Xg_<;[)]Ea2L08DMK>)+;KdWfZ>c2dZ[/-JGa=
a#@@/&=P_+]5Q:.Id36EX6+TdWC#fH0DYD,(6^7Oc,,[8-(5FC#J5DM,WN0T+.ee
9#RT95R5Veab8+=.C8W1D+KJc<d1XM8M10fJ3GFKNZ?@&5/-Zc_(8-)c)9Y[73=3
da7&T0,X8LA]/1B]OT-2.G]H?T]GXHKEI&ed\#.HVTX0(7356<8+^VH#\TF&BX6c
)6[#eOfSJZf/dLf.bfH(bPQ1VT_gAQ]0Y7XQdUVD-IA&3;HYLcVM5C2#UZd?N@;2
f7Y10;2>UK;0^PO\W<KM(@+JN@4T:V5c(\WdY+5,9+67<@=^8:)a?9CI-K)<4G:d
;IKL/9bF0OHC(K\KWSKH(I3N+[>_\^]+Z#>K(#4I>L<2=fZ3aHC6dG>P2X_63fC7
8F.A7W=HJaZf&f/0B]99GO(WKAgdG,Db+gOPMF>^EbN3cE/LF6a)#_ZJ)0T/gYfK
CRP(EUB+aKeFf)T8Q,>a,+.N;3B/L\0?_:ZbU>3B,-C@(g>6EbP=fS/GH[&gXD^7
8AEJ.7_A8N4PU6C@;Q^SX\3KT1@75<6QWP<#;_bb<b@/)P_YJFT&<=,T_bH7GC^0
VCN&C8=GIK>DWd;^YHF5A_@LV@Z&JYTK(2>KKLXU@eBC9GTOUEBf9g^bYC[+.QdV
^A\1.e/+T8OB,BM32.4dMU+4VSgZ(-X[F@D0[75bRU?O^Wg8.&CHR,_NQ56VVWUX
aFZDaCbd/:KUPH;8MEGBTQ.IS>3J5TV;f;<IMR;b48F8f,;P.=INgBbJd?Q5CGPG
<M+HC,XN1D(81;VU0V8O6]Y7ZcW39PX8Y>6/2)E7Y?)R@:=)8P7XPDO-R2aTL-Y+
CQO.1/(:f1?UOTT;0]032N7eS:Uc+=DF>1fb^Z--L8a)29N6::A25_L:JE,0ZCSX
VX_=Oc-JZR@XDV^2^;c63Q8689:CObJVE6PQYB]VDJY_-g2EY6FF6Q-cG4N@2K;S
^eP@FdTI+c_J2FMD^.UN2?ZcKeK4C1L]JDWM\_&>;^-g7KN/,>FZVb8Rc&^\/TLf
]9+0\0M8.(,F:8OaWNIM0UG<\Df;)&47KO76KAYeWg@e>db@4BgXX&4U?e^@XP8H
]5JVaa?&PVNZ\>7C)GIg:5dH(bG0\]UM=.e?A4bE=-<bQ?eS,5,A;>U]_[#?Z#R&
O2f3&R,T.@-Cb@41;BX):<#,43-J#@d40WVR)81J(;fRgB-g+=a7O<BR+IS1#)Z4
84L.D+]B<M0ZI@0[Ob0N6<2gc4-^:ETdJN>fcKRC[GUQ2>eZYBUE9-6=S^IZ1T9_
OD;?E(8e18e);X-&+J7._fH>JT-1G_L39^e&;_#G1->.8c:R8VUdAA5LQMFQ=d2+
_@0EG[M9A8;gA^?>K#JXB-6H0A866S\6DYUB4KB=R7&J9_BEUbg],_QC/:R[UZM,
;.LM,_OV5:SRPac#;Q/GJZQ8;dLLA4XR9f3CXKUBY6+GK#[Y(QDg>4PU:Fc8R]e)
)W9EgHd[S<3^G8(GB,>V1b._CD2X&ddH5@-/^/431_bX16SVKEL/CHBcCaC+#I#^
7HfY/^Uc+\M6,7f=bE:X;I@e1.]L[^S+,T^]B@d)1T+Eg\8LY5fL]B?5MI@+BP.W
AgcU4#H;AF7a.>2U,;I@DH#U0KN7ERD0W4g8SLQ#/L<Z]FU9URH#U3H67<b^cZ;Z
H2[8Za._M5bLI;K]1;[;Ib_:(C:G\:3GPb]aOC+Nd53H#2_0+Gc<(GJ@L711FVH@
XTHN<_)H,UEJFeSC<7]&/Z1:ZYU2K\^RAQ-0V\9\7eI4b55/@caLP.LM-fS>Q:/S
a&d<dM-?;#XK[[T2X/;1URIL_:K^TWf<W]0RTL6]KU60<Lg#V;3.88209\O)af@V
<<5[,>PV@CXJ0GWU>d4QGQ^>B::IC:=PUD6<NZdfNY5I]---a(K9(@,9eJO406ZG
2@-c:gAC]/]NH@(OWF#=2QeZ+?CE\]MPNC8/GE5BID;,_RY0HZg#F&(&0&#I.DgG
:(CNR5P0#b)CO7G8Z14]TWT9,E^1H&G_c5=R&RKTPU#IR49C)S>#Fc=2:6=ZaZ0c
)?Bf?2<TTC>ccASBHc;#\KPHPF(0MeTKQ/)#JJ3IB(H0[//4HbGQ0cd>,413J>He
>D:YBe=b)fOa<\L6)AE7He)F8ZN^&B3;R+(M9E0Y2G_Aa/8LP,L8G7>GV-JHb6VV
&5D?fZC,0&^RK9f6dgMH3:aE</D1E^OVFCbJFM/^]-\A4<aaIY.=\U?B-&;g,LC/
6:beG6_:f2TXOCBS)?H:LIA<EdF_.&VP69H#><Y7,>J0gLK3J7^QQ(YSBgNZH.cc
^U3b\-;a&2AW83e&V\+N5@8ZTE_VIZ?;E)3bQZ__dVQLa.Ncd_L)\)->bGJKCU2g
O<M?<aV=3]F/0R3a^REVO)A[SSF]-,/QTGZ[a(]LdaTK0>BGDbYPSI9FO86b_3:#
.Z5g?+BB-<;H=@T@M<?\_PNZf_\eTHaNaIL(a]S]KF>I^;K4Z?ZCEg3K6^-)(V1T
_ZWAY9/e[GL<T&/(@cIc]<&8XF1C_N0bB(AZ]8)_eYaK//BL).+C_9A:@]\QC>O]
:IHD)_Q[39:g&#W8KD+TC5IX9e?@TF/5_FMUd[&.IU0d:N,[HY]c(4a@cdR(gDV+
gOD_F^C=?RTa61]@/0MZf,\4[CFF)7d33Wc:?,SS4>5NA)Xe80ELI-e-L)aZLIO)
^IA1d,>]#IQNU_bUf-70Gf/Y@-FD&C#6DWL5:,<@Y-TI97>5I,?,/R(:g:Vf14D4
]5;0bJN_E5>,VQK\OfA8PB&K]MLeF\f&gG+^BLUPV^NLM9.)[#)7EX:XZCV06AB]
STIeP0J-89)N\EE/9C+LR\(TQ1g[((OZSV9-W=KWX><B9S/:=3O<SD/a(f6Q-Q5>
&3EfC;)D1+TbJ-CMGF>dMGYZYGD4^,(]\?8O2e&U,[(Q27=.ee40^1AB_&QQeRRA
Q)d,I/ee_>[_Ed.\SU3E8I3#6fUYMB;-I(-;B8dad-4A+7PU@Y=+4&V+c1.IS6U+
H05./R7Y+R0I]E4/gO,W:I81-N@=:S0PTEO&^??=E+9+F)E?c.7WH8Z?H2;EeKA&
DWg\40X1C4cb/+1PdT/bLC/<B]9:+gG2E0g^K+_c,Bg([8\WV8&[F@]8(d;OFN;?
#X?+?g\.(.D6WEVTB+(40W8Y:HZ#),577C0AN:J9&;?TIKd&T@:R#+<C^)&_I444
K8@:g(bG^Fc\[,.5)1<J<5SP-\>8c_?E?;WK1FaEL^O8+BPUg)D.eL1D9JE,U(8;
(PaB6/37ge]JSOIDKYQ/bcN\/,XIUI<N&Y#D<Q(.YE.X]L[SBbU+J+/06/[,C<)d
R3>.YcBOe94_>,E@a,A.)JgJ][3GMKI/WaCICFWg,9dCDd)bJT#ZI1^+<2CCBJZC
@+QHQ/7B?UBIJQdT^3+GXNF></F/.MI(<LE52M[Q>b=V&3>;JT=57)>W<7-d6+Z1
He>];ZGHg.FXe39F;N6eWg/VCAcZ>+Q&@CJbZF-7PfCR@GFWcfY0,=.@@dO2?dI_
JM@B(VbPZA;,BMHOY;=,aCM;?4F<E_8<,LdC:(0[Y7b=S:L[]6VVEA9-8DVLdT>:
T.efbLQ1U]TZ,TcSeg-[^J8Gf^;9E(V0(12B,bUg8P7(c<RPOC)BTa][0?d88[\[
(^0U[W]WE-URP\dG_^7,SK9A)Pe]NEU?5=XLJ@U)5[MOQ6[5((eB3IV=(RFJH3B^
?23>L]B&M9BP)ga+CcFY/;QHMA.1XH]bOD,G4>LF=FOcBB/[,gY<Qa(&WB8#gX9B
]?DJLBPM=R4#U19Ge::OgS,ceJSWebPX5S,\/[gK@967eWNHSIZE.32S\2[:S7e&
I_/:?F,W/&HU44(B;MTQ3I,?bUd(VOb?0C?,2cb8C_Ha^5cQ(BY>(#YfVKcI=fTe
_1fXT_W3),BKUa7G9e61W[CFb[,CEO,X4&?KJK<D1_]NS7NT?BAcJf<3&JB@PFN?
9&42Y_bZQD_+6c?HVX+]BP3PW7E&1?:8(&=I^R@Eg1OY1/,5D<A(82/R&X:)PCg-
N,Lg0+@Gc[MPDgQFcH0MEGJ/MgSG@;4VG4]=Ya/QFHQNVDfc[BGEW+Xc9?^:+_[(
=6<QKQ0SMU#YM4@=d>da[HJ?F_R;)/;^+EK=eK/T]V7KM<)#,1125D9?1BZ&S:KI
Db#X5:+PXL;+Y\N]FT7M/dX]TZVQ8^DX\(UC2a:d^XEAA@)FW]K.Y&+aB->2_XZg
PNFSS&1L^=J_53;KbLW\K+E(X_bf,.66d2gX4<K;G=aK+JGeXQT:3<a6N8^D;+cE
Rd1Q51Gg=ZTS.YJD)>&RWI598_[UW@Sc:].bO^XL5&SaR]++/Sbb\GQUN&YdF)+/
CU[=7O6.G;/66>g4>H0<3W=?2352JQ=D_TY1cb4OQH:[KJJ_\eKaV/WcBKB354/,
a^3A9>4F.H]B?G]+M]f;caILeFQg9(YI(C?@QFDZ/d/#;7VX0VZOECZR(HTbVLQ1
#We\dAOZ-ZHX[D^;2Z-]GC(P4c=@XDRTTOd=A&CH_Y6]SG<=]DM&cFdPP]9UEe4d
RHbQ_Me8(QcEM03)IK=/\0S75.X<04cN=ZF_)g>_2,2A8S4[1\K?]0a5M=-dc^A+
[+4=-ZJ5#)a.@8d.((Q=H9BP58;b0-:W;80_J7/@,TG<>ES+4J2]H/^VDf^U71,5
D8Y=UA19d@/P12g6gdBFW[Mg>?c.C2\5+9MPgFH7L(#ZX/G8NR,f8(,e1QdD[LX@
X,83Q^_13_YJTPO_AM9_6VC]bEZV)Ea4G1g0+[cEceHf<Mf.fJO/gL2?1XN4\Q8g
FA5,6+]CY0f@M]e#+QgJG]LfgUfWfcOb7H&RJ)WB<CC<^#Z?BR+dNSAGO8<R(4d=
E)IPI?49@dEBYIF/c2BB;>(ES+>=@H3SF7R#b4#D^H6O6;/8gA>BU;Gc[c(\e@4B
Z4[K.>RPR<6T?<FJ^,[;7+XHBZ;5<;E9E7Y^][E[W+VXT051NFJ5^]EcVXdX6WU\
)f[\>=XB6/:ReV:d6H5>H]3_2PX^#H4,^XO=\&N-TcZ.2(_36V\[.0]cc+c--9cC
MY^.L52MfIWG(JH7cg+-5V=#(#[<@H<VgTKMM_>UIMce-@\GfcZ>3R+TW9\92[)W
dcJ=C_+X.W<L)0-gedU;M[LT?0f(^\O@D82GZZ_=C=I3MV5[IFU=aK?aM@f.bgIV
J&90@DR\87)?e]J,5IRd0=/#_gdH9-RdSPbaO;EPLXa,.2-W:?J];+\,-VVS_]65
?T99==gNUL.Y@\],C#c[&8?OIQ4+E/I,4=NSbC)O,d6R+,3B<]K/V&[@fN5@RJaR
?\H,_3(PbSC+F,E,gf?>ICQ7CeJ=45?^??F3Uc>F0PY_:]E9f:P7-4TU7&8A4-TB
c^7?bA[dR1;4eGS=A.g>9d<,_gS=56g(#Tc#+Gd2J3IR9I5PX)QP^?DCU(.?<.EN
[1#^()UP-/&FT2a(M^)A)R2/d^F064885EYKW5_MQ2Q^]1FNOe:H,SS]g+-H5SI0
-RZUNCcg8@+TBU-KX/K#5bQ@7MBBM)5Fd.cJN5R+9=3JO4-4D0;\+eYSFGCf8]<G
Q4<+DD0_VM0QM\XE@7/&W0J0MBU7>I8&<C@]9H;&e)GIAEK8YDNc;R6AO/gJ2b\1
QHI=T=9<]9#65I#J;U,B[R\?B)aPC-#DeP:UI>763#AH=Qc08:I<ef<-\Ee(ddIY
,&TTbQeeX&?#F;B]\&@N1A93>MXK+>U2<.14SA>(LF1^Tf_YOJZ\W:1cb#=WSXeN
,7-O(0\W(;BPdKR9)>^Wd])TbZC;2RC5f]ebd[(RAJP?Ub>IGG9X>)^6gB6#f>+H
-L0dA]#Q@;1#_f6#?ag+7WGQWLA4A=2[[NDLN5\E\DR-?M1M,+6\-#?G3g85b;dc
?+EVabJb3?:c)d.CKN#9P),X/S<(8DT^Z/LR:&)8CX9/LY,CJe/0_VS?6?a:6I(V
<P0;Gb?Tg[XDa=5Q0?e4]/a69>]T7^0a\4U3N=HB;)^<:B5LX@F6bVX3>QP7Fa<B
[,&F,47&:<g>XVPQ-_5gIdTTb>P\WJ>bZST-UGaUc_8]HV>5C^7DL)[-dE3gC-.X
^FND0V5<Je;XE900fPJ)S^U#Z/5Ab70EE[[H#73YSCf\(#;TbRH4=AbcW@Q3#AT]
)Rf/6030/;X5ba7:Yb3F@:#WX0\-,L#8?1B>L&C:59#HSSDYA\B_W]<EAWPM+H2U
&:2DgE[S#+aQBY)Ka&K&;6g3#e3+=IKX\@P]O./XMKBP#e3?NSU-6Q2DJ@aZ(8e#
D>(._0KVJOUcLb79D:b#:++T?[ZE[MAIccUR>2EQ9MDMR>aMea[cN00;[0NG,-d-
J:UJ3L(a?Y;?HSHANcR#,<FKAAIee-0dBS\QU(g#)5d^_-fL?6(Bg-YO^8\\N\65
(1S?CMFQ\7#]VLI_?V]\f99;A/;e[:B5M^_[#)8+14fc3O\[ddM>PKdX_T[a)I)&
TAMZd)Se_CWS]3UFgQ8_SF(7QNSD&K-YQ@P+GW7OE,c?.HFff@B5:]:EM-8D/#;I
e<N9A^,>Y[d7QW98WRA;2@6(J/\caA^d[[F9B,===<,;fZ8bY=:O=a,8HT8.4MTW
Y0X[AaeK__NK\\AOAgO9IW<&1aeO9e3H&-YD?25Wf[(aG8e@Z9ecNdbU:59U3.PT
494A;V^@/^g:>+@F8e15IKPC)=O+G#KHLEa43RPU,fFRf&8aR\]9bcd<XecT/_/K
YO-QWQ_BSfb2EdRR.8JG2(OfQ8QN5#+N^]0-)Fb-?b/S^H&AYQ\dac#eLN:gF?-K
=^&RBYA6_B2eQPNe\3:>Z0MQeMI4eA9[P\88L(:?gC8T<7-<T9V+)-S?-4_9XcYM
&OJf=)WW<;M:I.?]g)9f-&M2AQ>&Ig336<3]KMcF];dbKTdZSXC<&[X-IgU08@K^
dg];@9BaS=+gcF)YOcZ)2CPD9/],3VPYa^c@@W)5S_M)1)/_GV)_IT3#Cga[N:2L
;Ic#a]<[-e193?W72?QMR>E?[Cf3+c]5UX0ZSKYB-b:\a05f)J8@?bEgCV<c.L.W
cdLIJfWAR3#+=\1cTf[aK/6>L/#>U#Q_?3NU9L?BJS1(]OI&YDY_9#gV0:a&Ya-[
e4E^9VH6@)Bcg7L;+T14B;J85FGJG[eTWJ@[Q0>^PW6#ge=O++(/&Qg3VO,GF#Oa
-3JP1)HbL,5E#/R-^1U<Qc2g8](7)]_A;PLE]>3<9g:U6OfW,VSGP^G4UK<5AKf@
S4AUDQ3(^,^I?5[4F.I&5-bdU26H\ZZK0a0a5H]#S>S#I-##dfJA&1.?\bda5823
&B:6N?MG(=,Ie)L_.CYb]+EN_5ZeH4da5T1R.b9L=;PV=<EG-CUed=aIT)S9BPb?
1LEVKF>(5-#,f7X0<,K8JeAPdA[5V\KS[O426F2\DgU[@@>-TUZ-D(Sg,VN-?W-6
9/8R6aFILH8&cPS-\;9#,1XC,(0BY1#YICZf2DD)Q.L^\3BM&>W4T)Z14\d@Z2]d
.XQI>)T)F<7-7&>&J4TAR_C-UaCTL+ff8YJ-0f,@PHKV]/=[K,8]=LJFVb(T/M+b
1//;T]G0g@C^S>+eE&Q8]PgL[fAeK,QG[TCgIVXS++-BI&D8DY3eP:f04Q4C8G8^
7GfX,)@^)a,622VP.N7<&&]1)+HA:M1.Q&VW:LN<N-5C9.+ZD#RRM8@FXYVZX;MQ
Yf2JVb>dQdN^:9F6K2d=G6SX(6]B=fUX]_)W:G\4X38YZI)8a1FX,JAM+NbLB)ND
\J#F05>]N)(1Z697+c,HFbJY&TI#FDbJKW=E<.c\,OODUXC;X9;VI+>@dM=,/JHf
,AE80V_F1Nc2]1;K0G+:\V.N0N@LAIU5JLPGOW:gQdJ@6H)VQY0CUVgKW]P3BB^C
QL_CZI9V4R6ZK)gS4<6P6b)ZJ1M/Dc4?ZCHEYc3NHTa.54PUE?>b\_=C)^C6BI-f
&-,VN1;-C]d8d6SVAb8/3.9@E@W\4C;MdACFWWQ.RTB#XTOff&1dA;P,QQ&R8)?=
AXUQWU(BJe>gb,GE>)[<,,SKRFcDEd3T@7;YaS2_W>GCI.<CGa.QUAO+DWG(#]Ye
DDZ7IY74LAL4&8GD;JCGM(72g+.&e__Z1]f4^][N1ILZV3NG5>7U4L)?[Q/2@+>2
M8WgBKVULgW(MR39fgQ81CbH,e[e#U3JHYgdRB6D4104R0GK-?2]X2Z22-Q86=Q?
f?/4e/ffZUOEaVJQDT[/S]&8GM9G^0C<eG;7CcdW\b\OZBTVOcXTX@c\F-)b::+>
CI?b1S_+)=WIK9I/7a/WII#KWgUXFI4\N9eZg3D-ed49@O+)<Y?_2)S2H0OD;bX&
Z(=1b8BLc?:;A7)R3N2O6[KPHWLdC8J:Mc^D?^K5T<ET1^7IFf50Z-1L;9^L)7c=
Ib](0O5QaECa@f=PV7Nagb-,C7HVbFTD2&X(]6Q1cf\-.S(UA/<C98Rg.E2D?;=V
M<&D6f.Z;T=aGebQ0C0J?0;e6DL/dNM<2Jc7fd:/0DfY<g4/8(SUReW1R[K3R=(9
Ig[IP2;S9XGRM8?UQ-+#BWaG][8bLP#RMO=d[_b5(5K+OR8I/\(Z@1\WI\SQF\-J
-[E7097W8?]>Ia=UT2JD::;>PXUE+W0WZ?#@RaZ_5+/^H,LOc+-Y^:D(,(F9(Ea+
OFJfH=,bXD0SZ9D[4Ug\R&SLY0E+W#7N/-A79()b?G1Y;aXe=(a[#;G0P11]VSD8
X.C?YVCfL_2(VSC@d,);5:?,9H/T,CQ8)FHE:[-RbLa:(cCb@AW:b0@P4Na6c=35
aN3U-556dE,WLQ(2YDIe,)4T@?VJC@@Te@bW-McV\(0\&aS]/0MPeH4<f84efVUC
_9gP=DN<HLR:edN)P>#P&L+WU[H2f<;Z-@PW>GS5DGfW8HCVC4]]QZ==JBec,X]D
:;6JNdJ+:@&5KT07g)]&_>/d<dE6eZaWa_a<b6f4B0:M_,a;3/4c^P2;S#8(Q#DT
G\gaDQ)WC7FV]/04La&A9^Y@OK7F)BLfB<e5RW4fJO(8>H]/dQ40E54SV=<1YZ9Z
+7(^NEEcBT/?FBKC^@WR02DZ@),N:=-aG>.HF.?#RbNeZC==M51c;RR\K(cg5aUU
a&>NWb?c,USGP=T+/<:1b+V+eMMRK0Va9^L(@NFN#dSV47gG]7S.0-(YDa(CRe:[
N^&9)-M>TNC37@;PN7+]g0?Lc&K^V>\c/.&^ZM.ASCI:^fL.5SeLeV4NHSI,@cH<
\X&KKL>3DKR.,_#.+V7eKLW4&cRW0>@^=O<c<HNXJ<XdcKE5&RPWK63.R/^\CYV5
_LUSX(3UQW#\[P7^g0BDMT:?Ke2X2)^53P9Q+dY>U1J8]WDX<GfV/5bQb.e#0SDI
2?QR@b6PP?QK@@f1b;C6<;3>)<_BBWdW@+D=7#X1LPVYRLS=U1A=IggQC4&.J9]A
?b^.W-/^eNRR^f&7&8>/AXXP0@_fE&]LaGLId9<9bf?8LQ6@5cF\@80PN=D:-<90
1L8.77E/8JZT,dNM<EfVZV;<J1b8:;V=5LG.2RT85K[2,)N/?VUUdQH&^=aJN&_4
3VY^#;fK7dDH5OCFdg)UaN0LDQNBQCeKK=MX,WU\d?-P:5O8S(c+5cB:-/\1)A?-
FN:TEFKg//D&EC+?/g_e6.dZ]bOF:?LUT<XIVZW.dBWH9[ME]0B=>119IARFe3-1
A#BA]O/c.\#,^JNRLB[0>TAW4VIWM&JL[JC\O<JMC\=7)GE,#1;IHZNKe+1_ZA@[
.9&Hb8g32<E7C4XAK7]c,XV<+=Y/]686VJH=-RG[Q8[7+64\DVQC4P+V-5-:5cGF
efedQNTcg>c7JbU&RHUX;NgQX0YE^DcTRb;0)M-bC,fdG-#PF#D2]>:/T]XFD2aT
1LI-1@Q,<RISQ#HT,a2\#7ff9eTE/;;K^HL+T,K1;^AXB?6RULX1d?QHVP.22@.>
L[9X:D#G&[=9F?eW:L6]DZ:6^^dVB\T26cM\e6,8PHXCC]U?70^GA@EWAH?SCJZ?
,LD7A@]Q)GX9EaB5O=7<KHPS;XJ#EIY@43.HCFTISCL9cQTGW9K5#ST=QT/HW8F<
[O1DeU8@O0/WMfAK7@,^ILg=(##\#;1MDL>g8d&025MQDXPA?MHe#b2Z19E@O]2Z
N9N2&cK@RI>_=IReW.d&A45S^?TXMK)RQ]HH-X=O)d[D&P1XF>;[9C;H#)9bOb@B
=3f_WW<0SGX;WONAJ\EY#]A,/_?N)gTH5c3?NOAJ\/IPM8b9F1TC5;DOSQD<,4]Q
Fdc[.5Bc1MEY6<JUIRJ2@UP+6Sc>8F\CeZ5B&,5_/g9ZSF=2EbJ;JS[]#N]./R4W
99b(QWD&>NdY5M1YO__f(#ZaK72cc+:ZALcS3Rc-UQV=,]42b5FCfS?VA&0WGf9e
_KQG=D=d(S_P+C)ZP5^C3TKNJH5/T5I3+N</F)0f0DgUDR>AaR46IM+:7:D&&Z7e
)@OY7]^SG42:M2M+Rd9b4-d18GT.QB-2?DEJe/7)[-LfV876XKFC,,8+IB)MX;gO
aB5Q/,I&2c,JeeD#VCUKLaI\Ic:,C=/@&I;YC,-AGX;fC?<@SDb1KKWO\f,4ML8V
Vab>4WJc_5[\gdGc_;J=IVFT7Y,ZB&W6-D)e]@))&C0+]6dO:K[RXMCd(,NL&FbU
;F]^S14gO)K[&OMD-aJ>8,@_\U&()&[IEQ&,=Ad96Hc(9]1?Q4geT>8I+?KUaJ=/
EHFBdYPC^4N61OBKaW6\Q2)WAYO[7,JZ(,R+IE+NJb&g\0SESOX5b=d[3_JV@9d/
f3SO8E#\Pb><E[XJ8L1D&(b^)J2JV942OR<;542A..MH-.f<]JXW+:M]&bc91/F)
Y=-;LMQ97#H<<09NeG3gV>SUf@UDVP5^^Xe1]FYA9#Q4#f:8;-XKgb30CF0Pc_GU
/VFe6[E\GK;)GORUZ.JBC>GW9fbBKc?/_6Pe]&Z]PP@Y+=ac&-5#D3fVBgIR\6:1
b(QD2FDe5C2UC_V6H20,]K+TagbN4W_44MEENR&YF^L_G78_,2.JARd0U&fQXQg(
:7Q:F\O1&cYG_^\A42A,3S:O9A0(]bDT-,WIRSKAB(FPLZZSMZ?S7I\R.R]3[X9b
:5@ISUVNTD_[N5c0d-S8??,@29BFG1^11-f)MgQ42O\[WKC/<3]WEUUJY?TGS1ff
7Z/.A>&76)S?\e5@d3IT>L75(+1=)AW\7e,M(3)1#3?1dVgeOTgFC5^S;3&XeT=1
bf^dYDaKJc4(61RC.FdSac;&K8=AUW\^G(1-7geJFR\F3(3O=;Y9UE/QOH=8&9_K
[3#KN6<eYW\#/@WVUZ5[HX3+3WLO[1T#&DQ7T4\:CB&BVAFOMbf1c(@,9DT]F&(a
C&#)HBc4-Q=8W0I8F:#KTV.0ZF.,@1-d+CAd0eDb[-FbN(J+Q8&,1O=S6a76H6eL
G1YN2S8V[79-^S<1IL:/aZeTBcZ3J&C9Mg4)gK.&L^4?KC:S]X<[#,)V9@EIMR_X
MHN+:?b-0b68M,P-?BcT.B3#eS#_:)C.)=&P>9&3;-;>10X8eTEA@O8C9R?WO1WF
X&M;5T/E5cER1T,_=Q,/J2374P_F1T<-M:S?g-9:=U(8DLA1]H)3Sd;M232ZKGNB
cCeR98Cdd.5YS&XJ/fb09F\5&.:a(LN9.>&F(&9\Kf#R;OVUB]L_2KE#TW\OSW-T
[FJ=B]CJ#D7(.I&WYWBbc,A76=bT1;O>Qc0C?N^UB[:E,OD#Q9BHdCdGC&^O6DeZ
@MVHa&Q@A4WEWBd2&cNgZ0ZdKFISD4Y1629d<7S3b@:JcSA&JNAHU@>L5K@0aXZS
N6@P=Da?E47E^GDS3-L0\>[[IUT[,57./,B\A#7:H:.6CL)2L29]g9K39M1WL1HA
T4LNC_P]N?W)^f-C>BA=Z:D6f.JZ46;R^VgMI:>aFZ9,/\<O4g9B^44U[P/94^d]
J4M@dM36R,\XG)+QKAIJL(e-ULX6)+a1eP)eId?,J4/gV[c#gX72<?FE7dQ_b(LN
JbLSG,563<KG3@J86XI5&V4,Q@YHBMG?B@\&.@^AeG[1^.;/\44#(HgQ8#QT0Z4S
DdAGc?1gGS_M?:9(VTJVDLECV=[ERFU(O+3WV2_6TLA7<JA73dYA1W,-3XgW#,XY
afg#_U[;[R-8O^HLFR]W.Hc66GV[K_3R:JRN_bT,F=]AD>^Meg@ZAYO032f./ZRX
;RD&@F]a9P/:a=YK#HAPRK+YIKFHU@ZE(J[W0;e<NUgJQ=)3BK38^V4XGMYWgX:^
6TFHHX@/H,XYV67WT@1O1M30WGQb&<3G:+_g\.?[Ygd=3.?#JF]gAW>:#YP4W\d,
E#a4F:cG0\FAME55HK<4+OP6Z/C++KEHe+NX7#L]0#:dH(BaSA6FO0>3J\_RG1-N
0JDWP04ZL.]U^@3/Q^gG:XN3]8Wf(AKSNeLe@#-S48\d)SZ=O?B9(eH\8[ZQ5@eC
2g(dBT)J<3<;#H=.^[1:N)2dFNM=Kf]3@#Z+6W5_&_B(&KCFZ6ZO(QZcb:<b-GX>
Q/AfJ@g9>9cGZB^a&.X;2TJVK]Z/+.Z#=B^]BV^U-S1FWWfAAc\eJIW<\aY@K==[
TKa7XQK:IA+=.e.=>((_Nc4[9O6.U01F9.-U#7=bF[Q?N.Q6Kg6M?MG1e@4K.NdH
6MA3=.T2F513GD.V;<g]QP@G^@APWWHVX2Y:#40B4EVY>5<(.-6a#c94NI/_-dg^
T.6Fe4CH3P_@UD_0@-3CGT=PfY)Q;<R)LR>ES-L:LPBIIc6/Y+Q?W)&?UAC\PT<@
RJX?DFKVM+R-8=_8R5.&CFFYU4G),-#YDARZ/.,B\(>4#\+&UZYD_#JEE,X\b27,
D[:J,GEY+J0;=Z>V8#S&a\.Ta1,KC0S0=&e<d_7d3b7771,CE&/cX/+Z[>W=bYT4
)c9W5J.)M;G/\8e7W;HY[fU(Z._HeA#4KFK#UW:5.ZV#9N_FUZK:\+O(\I6>L0>b
H(Ge2@RY6?/bVPKbg#1SA2,[Q-)2,3OfT@U4ON^B@D=Md7X&[+8OAIQ^4_R.;,R7
Z1P3X>JM^@Q2:H<=(A=D=EO68\dQ1M/)\9f36(BgKZ88&8\RG:a0JE?+#IaD_Mca
)R,<C-15Rg44)Ta.B2PS6X7d@gF3UPMD:\+d#FU^81Y\F^/BPU=;G#E/Z;VVe7Q:
g2]A_2L)XQZ+XG:C46[acF2O<>eU/<gc\I94_FG-L?1CJgN1<bgXQQI_S^If_[X;
cb#./3M?097\T<IfRG_,8a9^C=@L?>7]@a,G3AGHD/91<1HCg?9e9&N</ef?M5F,
BK9S0WHNaAeF3,c#S_dRL=TRfNM-d0bH9J1@b846KFYSR9AD.Y\7V3156,=c;Y;?
Z3DDJGcbf?1K2T:03Z;<QM70=J.T@+:OW+WdfZ2N4GJ)A/E-9159+J78d[OUL-U^
27OGX5e.D^JH9C?c>H:VVa?LXI:<4Y^9U3XXW\fM4)a)_&I@<D>AKZILK1GZ2SCG
H)+V3-a)1/TU5(V?/\XZcIeC+Q0f[0d3N+A:UL3>&)QRQ&SV@T1V>Cd.VLC4gW9H
2Lc[-#WQ[Y^+^7SK]E3^g<<YETLECb1UHI:8\&Jd\B;94NJUZF0W6?05Fc_2,LO?
#9A8:H9&R7]#5<9Yb_V5Ta1BV23N[c#I4\@(_]9>AYQ\04bQcfe(1=LT.WR&PQD_
4\^NOLZI0]P0?_e8bbGX@Y@U6:7JEF^#Id2KM_8[NSVc0Q-Yd,WR-7REI<7&R;MQ
TOgN4XYd0_.2V>S_16:I[\LHGLC]1]IJH9d@A-88.]1fg:;GA[8GB<N<+6A&8NP)
0DLP.I0&8H7XCYJ:X7N(HG#AdK-U]O2=.S>\W--SM\Lc9=_00FO,e=<2(MA/8f_E
W&<34VV8EAa3SV[b)3J(,Q_FG:[=4:RO[R/.#N?SW:64OK,SJT1bBHFgDZBXU5:\
<10<(^e_,D25C0OeeNO32EGG\80SSC8@bc2c^\IdeAAAIc,;___G4A?\33gR)?]E
UIUbC7fa?N5\N[/4dddg+:T0ObDcXdA=4<R6SfBO+3V.OBDFcI_/>.=TQLfW\YL2
BJPC>c0fYTFZH>M4O66C.g-1__W=+I#]O<ZW[89LPP9EW)H=6VB0e>^IE6H1SZRb
B)Wa7,[<U&b;1B>HMVO(::RLD2&M@<H3SPIJB3(AU,/7I;M,_O[O/J[8,T-0&F8P
CGS:M-.7+9c[7W)^11gB\Pg0Q/F,JH&gZ&b=N@4\XZ6:,ZVE/FU#\_.1#[4/:+)]
2_G(U9AB>5OHR)-QJ?/_c6JB&ggG5[LDXY5MEL;WfA]2_3VGEb+>.;..YRa\_H_I
8?KCG5;R(/VWbBgaZ6H5W.38F@YGC0R<aXA4&+W8X[46dSRC,YG&DGeHEL><bU#2
5/OEf=?cC_)c/);ME/4?2M/4\BMI=I_(4bK=bae_;-&JcL4=,^E_XR8_.D=(IG2)
L#2AA:BO<=)/\^M?BQS1U1L2V/^a,B][N3R:+9.7;),60XOaD8X;c@Y_bbQ[7:F2
E6N&dc>OLULGM5H^FSb/1:7J<=GISY4W[?aD2P^ANL@NKX[:1#:VPL1^,^SW8U(D
72RY<bgY#[V#YP<^N.SC/0:S<e?FVK_/bg_3Z+L2e#(Ae0aAWNVAJ5T[B(8:0/)=
&T^@JFYdEX;4Mb[Ie=RL#818;UC]A]@Nca?W_Ja,FC/XVcA@\Q/MV:S^VdULJRe9
6(9OT?(,#=g_#7(KPY<(DJ5&cGGO@:2;Mb<DR])faeE:7BGYa.H]3NI6&dVL.<<L
R3CZ-L#Rg,[&KVSXZK:Q/0;BA(1P^Q>[&87(<COJaeP8^R?0R5^@W;JKCTO1/G1C
g]DT#Z[1[<LCYfS(ReC_a:T#U-FT39E:H-BU\)S/\ZG(UHe3QQ11W8PN-8CfH7L[
V&g/,3V>EbE;ON@=[JM/g?PSfb(H^?VZJ.fZL)U[-64BE<,Fd4RX8WDTL8c[&),;
A;R>;CPLMUK7(VBW4a8bNH3NSD\K2cRH.XaS:6HCY++60c-V:,Y_e0?N[[R=BYeU
OSVe0Y^,/6@<#cOg_^^I.K/BIf[bV0(BE<AO=4d+/A;U]7U>81:?Rd&13OB.;3S_
>2ZFG9a);:eW-#;08NI.0@0VA>#V8RW;1EV@L,V(Q4>^0A)0O62QWD,c04,@@R(&
/7ET@d11&FS>QJ0@(dd7Y-e;?8GFU_N4/?RLEJ5W?Q[eXJ@>c12dM]]eH1,A1LVg
,3#>g6&@PXO@eK_8YUS5&7],.OY6TT2aIa0>?]J1<9&9Q;04QB>cCIUX/K_A(5TK
--8NA4_Y/DRO_HQ9PISG,8YCQ.^E++8MU?>f:SC\/>;D-Z&J27#)A:;@GGH]@:-R
=/G=g4T.5KP60]S>GcKB[]6e.45LNOV[Y^_G^T=]gM+>(11_bEJ1EcEQ[R9C_]9:
.:9e@a:_#M?JBUJ8>]9#gLaHd))?^<TWfPSKEBVJg)?S3;a)cNV81].G2=ED_F-6
KBCE++D#Z_SXQS/+c42gI.dfe.V>B5eb&65.MLY##X,=#C/6Z:;0=Gf623FC[Z?7
4dH_./_927Ye3;TC>E;b6C#1L0KM^]_5@f>BAFeWLABfd5X+YD,F>C2gQIa(NJ_G
e48b.Ng5JZTCOORJNe,/U01;HB4:KTP7[;3;>RQPPfe1M:LbbYY_WN1N;B7Z2B[=
/SL\S=9<#SR3S)g_N760e-03fUW=MX=9Xb@O2;OQFE=/0GI9.-W1Q#<#I8&PJ45/
Bf;/fH:PSW+RgcY,f];VggNJAg/7T4M8>#gPa;;0H+W6dZU88Xf10J7^M=dIQ#2A
2bDbOAJ?S#JO]7/D4J43ZNT9b4Z-aObP4_)@@GTDW)OR9cOQ0Q6A-/Q@Sb]S(7:K
\.OLbaZJL9AP):8(CEeIN#XDc4J.5E\QdgSWQ2,JcP2T;DfBO=DV4B@_Ob/;GSf\
OH#X)aVP,_F8F7_FDaI=FM-db,Y#5<FR)F+?d+7e.:1=LL.33T(9eE4>8cFP_ET4
R=RQ7-SMX;CHJc4(0#f>5BI726(W\fMPc0NHSJQ^R@T-7;313:W/,Y]SM6cUG\)B
X#-(e;Cd3W_XfTR>,^gCMNU8-fFScgcVV91&=NQ24eIV]PBHa/VSc=Pc/a@V)):#
RDG9cQaU^>E]FdW3N.5FBR/)NVKCAdd,Sf&3]0]T32MWB07-[;eM4H7#V)YF0gUX
NbQ5.F>97^cdP,Y@R&=9EfA&)>OCMLCc/NU[aUDeHe4UW27RGDV&a1a#6VO2bTb@
U8QU.;_gWS(/^gV\\AMFXF0E:+N7O4gV<K@;;1Q>H9=8:2C39CGb(.NUaNb&gJ9+
0aQ>0QCXaRK3<W<@+(X,FLfKY@QL--8AYZ8,S6<TcM<+2O1O[Ec43Q+B@\WcVbNA
[Y;7b.IL)]CXNJ4+\2]aT589ea<DFTb1DQI[Of4)Od<FJ)5[?NA3CB@B>\&P9b(.
YBV>=]H7#.I^Z/MTQfN).GD@+[SE^6IB=(8>(2?78HRBJ4E9J4gb:)HgWK?]dB:.
A]Ye#]5,6?Z5^Z=46+G5[4,d)Ta?/Y:I)R00OH5N3<+A[fBGeE9Y_cI0Y)K>gC.G
5HA13T?@VL@TTF0;?K+FO8[P&\>a#Z/@]cb29Z0JR#C0f@ADOI+_IO>VQ[0RAF(N
K>+JXFH5PF@2I;4I3aTI2DR(=A=3#X,_3:F6&G;d@(A.^:&K<MTRU?fZJ^gHdHAb
4+LH?]A,fe5Z#HdVT1;2g&c<-;W]]J8?ESb\XLPGO21(W:bLbaZg#\G6B[?UaN6#
dS,[9Y+-DLe[K@&U7bFXK2f,F-gGE55IKacaI9(>8+6)-TR)dS(#NAYW_G,d6MKf
-R@S.G#SEZ5@1D2I3:@-VXT^X>SM5B-TdM,-#1MaB;<-ID<T[OdQ#E^Z_e0CWNZe
R4IQS0bXDI7\:2aedB9eCbWV^L^c]fV<B:^(STXTT\Ef4C82>X]3UIN^bBRDbCKE
WWdR2>3^/IQe;f061Q2.d,XY\3870X\=15C1&YWR?77^@W0QG;Z^REfOSY;-N:6T
Jf&0WDO\,R_Y6HJ4/XBUT1f[GR/,+?+EZW+3WgAY>0WX=,f;C5L6KaFCXM3d2RJg
A;Z,Y5\.f53Z[=ZTgIW)?&@/U6]G+dBC.6\ZVe&C54ZUHGcC6<7&1bM90;J2:F(?
UV^G]Y[24W2&<PWM(\TD.O0,CXa=AD:YT#GV#9[e3KN0?73.P>=2Z/+></^97^.>
+O]LdZ3ZD4K)Nf[ALT/ce7L:A/LFW/=8).:9FBRaD4>SKSg][IT)]/Ae?RT/BX6g
aQdbYW4\)KK8<(Z[I/W:?6V,7dWD:(Cb#4V=EXR]FY#.9c[aA/&XV7=dQ(&Qe:/7
P\8gBSY?4XEB@^/834/0U31J;BI).Q;MBG,,HK5CR>@LDV,a_N</PD@2&/UTgY99
Jc<M,L)]].HFKc_&JT:63JZ#EV,I&2-:K2&cd[DKG8JETF0>Rdb=7^R2:S5[]Z2.
RVQR(;;<JH(J.V5cV/4PF(TSe-AY[WVMA\[,FLE.,@D:P&C5P>)5+]1gI9.=6GQT
0^)4SKSJ7J<E522[UF?XME>e,_00W/;K0^aL;dV):;E4b/Og[ICB;=Oa^<;5?W(Z
e6D)+T<6MZC,HeFT_(e5(.V4CVd=gW/b+(27Q>9FAFN61D)2cFHDeXdH6-.dBSID
aVS[ad7\KCcP:XcFG+5JRW/(PR4ZceV_MYgIMDY=)UL238\64[O(XLU/UGIdgFS4
f4+X8N22fY4bN1;cW<[[CCg@XJLG)K_Q=,\1fR<f;(VNS:a:M)ET/TQ8I:?E76((
9YC\)+;DP<W_SYN)>c0^)X&4(U^;bE_<^OC0:=:T=HQV:YM=67G/1fWF,/,[9Fe)
;8(A14:A4+,1V[6COY#LG1ZSC[b7W2SaN#1f-A<_2?P67DRLD\NV2f@De#SccO]6
CW7#Ib#S#dE=N5=\W:A[3YOZI>[c-E;b0V<=E&J9CNAF--gXQGC3E_.D,Gf@\A<J
EbU\,NV()3BK:__b@/+P)F.AFJ/:V<eZ(VV6E2f?];b0BM(,0;TJ?3ZZ01HDfL5<
e62UB(2R)YHNYD,9+aI8\adMTaRQWE<:K(a?9f.:R\K:/KF)LCgB9,N;6QP.BD.:
CP[+KEE@)WWT;U7NAMXV;T)87NE]BF?._JX?Ib@LQ/Q7H<#e--aWS3IM1_:B?NbG
6/PRO?&9_.Rb3aNHNUc]65V>HWUG#F27dB;+E2a.NT)Ze>)c2-))HNe5)2EU\e.B
)I1)a?R+;-]14+)cOD5g<3]KV^Fc39;W-CT[-3H?aE[c.[)(TQ:bTWc&\D@ec9/K
@>GII&38I@:I)?X\gLQ=@g)ecHYY,.(P-<+^^/)b8:@EcO5\9&@_+:Z;QXb2LQMP
,,:WT8D5VT<9@QK@P&[AI,I^[89M2;;.]G/-S095E6E?[K\9LSWS8=502FeLB_;:
>d<+5U#eTce94I/c,U:TfW2,L&aUd:SC7H9W&,(^1[V+;cRD?&4,cc/(RF#M0GUY
/-TT\)4P3U:bL<6_S#WaL-gP??#1R@FL.-9XLYg5b/(738D],84=;c])2K_]^4B=
<\C5JTF(+@5K7)<V+I^Of(U9MRd3YREWWdeX:_OL=54D9dM(SD=JQ-f]CM5;8CKW
U^VV.(S^VH?6#O#DS\P6X-=].>2a@4\bgHF=VT?:Rab2K.7YGLHJK&b:f-W03B9T
Y:+_@&;=96&<\#\N2OLaSMbaRd>#;3/H#Z,R0eb6dQ&/T]7FSJ/HfR^]KJ&I/,CB
266IUWGAO+^5(35@CLE663+_I77e9G;c\BBcaPW8?B0d0cYbf0@0VDAA8d]ZS/0a
ET^]:^[F-K9&_3;V#6,Ug2Z?(G/1TD:DMc3G(DV5H2LZ]46.;Xd=(eF0(Q_cPTbY
IY1bW&<9ILVTeZ+J;bf8V2G=1,:7&5;(JEU7+)<((MNTQNaBHR6d.J\HRY22<DBE
PSOGH@K/HQ_7&PLE]I;HF-cg14S\>c;P4#C^F+>#H^g05b;XB92e#;2/,/[ENOZR
EVC+(=@J5a(VFb=U^6J48LZ>ePK8E;DLMQ\[\]H?Q(VN=J1gDZA;NKK-D-dcWQb;
I9&=Yg9EU3AHf<)FPZVe3#-a7V.[L@3UdV,6[=5]J=,Ya-9A42bNM-Ed:UUSJ]^>
81[ce&RDMeC/=@5DC-g69+]V5O];Ja\?c5U2<fZ&7^d29YfN&^2LN0(;#Vc4f0X6
[[5BD2E?6A1JfYS@K(#gcJA=:9AUcERFX3F)./aGG.Kf<MK&#E9/:5AP3K)bc[63
@N7@_.2c/?^8Y&b]45X+_4&#3TO,YfaST+\3?0eU?1c9YL\=H9=HgcbOWg:1N17)
5CILN+\DW\@/]7,Q6>2b]C8Y;_fV[@P&1G=7RMfJ+&-cFbQU2eY&S^a3Q4P5f/>#
DV34QIB,+>KN41F;A>[G=4]R@P4g@G?9M&->Q-J(Oe6I#M[,,&HTOSAOO8NHaVaM
HNACJ#UOb02\@=GAE\;[@:_EWAFT&#=eO^c7107L^#>@45d:[1=9(9Na5gTGf]BP
5PLVO^4O#K@Ma1aVHR;TW^KcHe6eA3AN&aW99#I5Wf?.^a3CL9:E^21S7S+346NE
-TYX7\LI5<c5J;31Cg(7VX/^&Y0X=:#-DP,G;<F(9J@<g2LF^e9_9)L.Hc?MB/]4
OMJ0P_AJg[Nc@T.@gOe]I,LIVWb-D:<beAW9\(1SbHJfT4#;N.0d]SR(d>DRI+W^
(@;A+M9_H^R.&]/?(B7R&<++TXOMAI-\=d-RDJ:=<fD<1VL]N2[P;8BW^W/PcX9<
_/(IKASWQe.W\Y:G1=6aJ/=/EJgMF8PJA[>eR&W<Y]B78XI6K<N\P^c3e-;EL,)Z
HLF-^SMA6?1OHL4R&@#Rc\^X]:8YYO=GN?(R,3,E3@A4GLXEFWSQNG\NT&M^5;B.
,7V+SW^/.K&L3T3.]/?e2^N>91JHFeLM:M/U&PASg>]K<CNN#XE+Na/TEc;b5VF1
)T<d&D+.;4\NE@D.e&3I;;XFS:,^1A#eL8ZB7WF#MAP8CCZ;[?[K^0[MB0WGTF9d
+g:dF&R9F;Z5PG/&,O0\RO^Z5VYf6]KdLKJ#5)XYXC=?&)9=W>gC&Q01c<,DI6XV
fOJ2I<;.YL]Gc,[@,OM9^N-fZV3P(Ea[#?IW]d/1CeE(/0:+O]&10b#;80>dgSNT
]d/86;[Taf9TI.,CAC7KaSbY>1K=3KOeFT;MGA]6IFbCbA-J5VOV?B#5D]:=3@G<
K7#YBC.F_&4g&1#HQ>X-g\CGK[dIA9L_HZbQNd\ccILWSFG>,3HC]@g]>WA:-Y;;
fTe5#X2&b3\dNA(ECQbSXH[dR=d<6GQOVTH=b.F/;(3OMf+g?P>a4@O:1@QN?_A/
VcUe/^:+d_eOdcY.<2f//)b\g_;AdcF^4BY6V#@IZY5/.RG][+A)P+D/Af?Y2Q^K
Rba?d&aTg4]bV110D#1EXUbYd?QD&&S#=1JZ7b03E<LRad=&+1H.:#YYV)#/XV(?
KP-YE+?bWaP9]]b)Q]T12KW?J1P=A(eYQ:<<GRSA17Q;8IdaE[-ANM^#)B7gSR<U
/6=_O0EQ1a0[N3M7Hg3dS5ZcGEE)Hb+#@/U?e&A_^HW_a2)7GC87N1J_:N2^UX)W
?b/6H3d7-0g<\A]J,K6We-/U3>&?T.+9=RZ&5:C0c@0^)#UZ&Vg-HQV0TC<#6OVL
J8c_eZFZEdg-b;&-.BGMKE;KJS@2<;[R:AgHE4C@Re.R\WO?Q\H5A4Z[X[OgB1Y\
8CZ<1J:.Z+[TYN+YfXGdMd.0;b;CfgLdI]:4D<91D-C9=76PO-A]145JS])bR.9_
F)IU\A+ZJ>P3J?U/K:=Jg[V\Z0-DR#)eBW-5A:A#Q[I(fg&U03FN.?RTQ]_:<X0J
5)Wg#&)f,c=K(Sb@1-(fCKfU>JFQ(+CF)e([-Ba>=+K2(+O=Cc5PM>+TRQ[f]Z[g
:H&Q=cLG(:Lc+3WK)D:,;_4aA1_cRF@G&-&gS/eT5UR_3g<81bD#P:1dfggRLKO4
]@GKG&QSX79THOA3^I);V1\e+Xb>-^R>O>Y#FQULNOd,A;4gQ/a&B>7@1VF4>&2c
+SM;;ESNJ0-fIe=S]e@P8ffM.=IBNQX)#(:e\0Y]c_B:VIJ9(ZL@I][_AB8Va_X1
E@EBE^cS;If#H1<DI,g(8JT.=;\A@WOC4H[+D<G>Rb3E3>fT@B4[bScf<VQ8P77]
VeN]MY;Ub9U4@\Z+9)gQ:?>^80L-EF76.BRd[39WN[G#/5_51[X\)^;Re54T(6ge
b(gb-5YXcT7a<QIUG::@B<A<g=+b,K80;@84fc?Cdd4\g#X)#ZL_aRa1YR:)=Y8-
XKd4==B.=Bg=D3_g;4Z=7\]+@4e]Y]2W+-,RZHU/79e3[K@#<)RFK3M_LH9Y+cKN
)JY4E.9T\eO;>ML2_+KVO[OPa[=HBgN8O_DMW>0H1[B=#IQ@1DG(9.+If14G&EC7
5,>DAa\7T8)BBd\YR1XLBP+cSDA@4IT222HF2SOLG464EU@+:g7XUD7HVIO0cF<^
V+EMG;.].)&AP9^Y7+O(5EK^67A_gI/?T;1V]#geRD?V.I2+OfH1^(E<070LFD1W
/,Z,WD9<Xd+JE;E4KZK(L9(P\B\SS&fJB\)/=4XY>24(LGb+S:aH;)gHXJg^?)YU
cE>N/I]9N?VL&,(&gU(;#,_7E27(a:46E5e<Y(1(6)RCI<(1Z[1&X7d^H/:<S.+6
?EYY\RBKRX[@5P:<-4S3YE9g\=U2b?XTLSMJL=C,QOPY[V#dO_DCf;[aD.#NG;^;
+ICWLIdC+>1AdE5B,b[^C.g22MCSMO+MdfGZBS>-(bO_-<M1P;f#.0T1_4CfYef<
g;+SU1?#AW)TPAe<aGT;7M@NH=8A35P/Z)]\Y2S>;A#GDV10\A?Q7]Y(]<KC#-]g
Yc818g\2@K?cgOb/gMRGN6I>8EAE>(Q^(Y4-;b(E\M?>?AKN(eLKM.V362(@GX4O
2&./?@:I,=O(fgI?WgX0aL6YT?FQ-X__C3d:M_c-_bXJA#Rd)HdTL8SDM^Q:?([E
&+Q-\(,O?Fb6=WW9>5+P?BbdOEIAa-L7660/Y-<3:\_D-)/a-:AF>bMWe1WKF>(L
d?Dd/WCH/R\QEg^N5=]X0IEHBJI^90Cd8UA^,<-UT8A;Q;1Fa9U,1OB_#KBX9EF@
5#F1c#]P9f@K_+6^:5/d)AKX(>fYJIe2P:eKbUP4e;+9U>.O8]bf=I-S5_?N&:-G
)]:d+aE-ILS+/4&A/1c/G?gOSPP0[Ua:e:@R/C?&Q/a?bf.9L2J?He\X>1,]X4C^
;^,P?174VgQXU<+CS077^I3[#N6PN4.7BR>cVMJTD5bd^PX3])+F(>g=\/EcJB/8
T?-GW+Q_Nc?b1-WNXZ6JXN^1WD7:TPNTS8S<I4Rf5U_14HX5F1K2H#1/7f?8O6B&
1:TQ+X6b4?_H)eKPAH0^)?2,TP2He>?3g[YBH;1g;]UaDC^6W2O5G.ZS7V[]?HE0
D-5X+F.e@8&IVXaOL(-0YC-QeEFUWC-9KYGRSMI&ddVC3NP-1]G@135?H,O\2]1?
ZcGg#R9ID0KdO[9(0cTV_2.@5-WQ+X3)b.KVIaBZ_@H,SeXP\TGU-7[8>4e-XN;]
RU)>KHb@WCK?gEL?&DDWH#6e?XFaLJM]K]=a[_Qe_G#-f?@&c325?_6c<\MV#_(W
[;#N-fgaW1UYS)8,XS2g-P?#8V)fPcK95F_d3Q4;S:/QK.Y-YbA:P?+#aZb=;4<>
F?Pfb>B4.+,R5_+V5VEFSZ?JMJCS0LfN4+\C^9d\0ZN>^d\TXQY;B1):/dDaGRBW
VH(@fTMSCLQMd?[T/MJ0g9];^e32?<<;L_7TT@<XOY-EPg&U2fXUN-b>\Z8AaHRg
YJgcBF@cL,O^=@ZLcS7?K;6eOWJG-OE(94T5<K:4\fINb>ISJcQV?V934H:C_7HW
#\?EY7:[7CFff9f?b0)Ig;ZL]VGf]15ITFC9gfW[/X8d\HW3/UM3YX9)J?6;2cNT
P]+fX#WJ>)7Y1P3CdMC<G)QfYcP4E&V9IVH]8R>8>VCf)<e8[A2Ta,JTE/OC[fUE
//[T:LB(B0K1^C-Xcg_UJX6_]PP)&>/-_4bP,U^g1;WEV+^H@EY6eb1,BZ52]-9O
7^Q/-dg#,^=AXLBI7<BK[<0dFf#.C/(=@d8B<>U:ANGYc)eP2S16Y_e/IFA1D_FJ
W&=Kd_?F?WCK],NEESe/4/GJL[V:@K^Ud4]Tgd[OWT5]7DQN(a=+V\)K;@aSgQ7K
R:VF59Y)W+aX6W//dH0faEWYF#O)4-]BVUYfA./8e:/JcB)8f[/J=J3&F\M>78eO
CQV6?CPSU96DC8Q/Jeb&#4_]\LS&9<OYa7cS;U:D0e3,F)V<KK8bH0PP47fH7OAC
GU,JO@Nd2J739Y(M/[G31TS8;(MW.^A\dA^KQ-V6/(dSfX=KeM-<+E[7VWI_FQ0K
8/VeccRV0YF6I.F(8&+;ATR^[Wc1M;77&U+e/45+EC6^9V,f&6YO:\:Y(gI]M,1/
:b_A_PP)(BOaU<Q?d]<6dC0.D15/.UHK3L>FO3a8D+>c@aPKec?gCSdM<JRDQGD5
@]\Lf12S+-OF2;g=?E:][IBSF(0I3OP7BBaNV10Y6N14?SO_CJC05#d4bM?-37:a
Wd:SINWAS,b3IbEG>#2G9;9#GSOYTV_7H6V)^[T(CZ0P\YTZgKBa=OZQ=f;FScS=
_&Qe1TZ3P;,ZBT8K#F(4<<:5cO.FE63B04C;_P<=323ZeXXf1AZ]\2S\aDLLY5c9
e:9FNSRH42\.L)P5>dKYAf1>VV^g7K^b(.(>_JU1UWX)NIg&OSZ;4Me[84CMT=_C
O3<cY_.Y65#Lc=NeCVA14GVcIE2V5Q_F(#4&8cJDgRAbG\)WQf>&;KE1_eUcURV;
FAMTM3Z39.[N73-WL_)d:-;E3Uc\K6:GNfYOE+HIUR:)0JFW02K3FW.9c=8,:UVL
Z=OD_OFNA\.ZORR1fM<WMbL?4<]KXMG:KM@QS\D)18?7S8\AbG8g005.PJ8D49]b
,AF,4>9>(4cHdgXN9/IGX2SQR5,[8\BQO/,0H_FB=)>Xb;QDO#Ceg20;5TbR0J0b
96/fP_eMWO0-OY0C)N&YBcZf&9B/6>)cR]3B4bK0^gCS#.2cJJTEe0Y;9-0R<VYD
J5FVN:J-eGWDR:Y.G8QNX3NY#J(EF,HM1^XI@Gd3JAg?1]7RBZ)^f._+1Hf0g&b[
;:6e;5fSXBLAdDLSaVBBZ@,#A;@7IO5(H+M>S(A+438Z[<?A#\36X<+IV#D+d:e>
TWX3#0[DN+31IN>b6:,TV[X7]NG>05Sd)5XM\0>></(6J#M3P@\#;dHcGMee9F\-
>.Z#AB.J\@-G#IW5(WQ<NMGA_9EQM\W\\Pcc.6>B115IQF@F>?Y@O\AV-ZA1b2_2
;?Sc,RE/(11\0d^#D9SGX/Z)TIeW,aaNgg5O;GB&^fR36\HW>Ob&#GSX?aK^OP]W
_^bG?O@6,MLFUcQW)Y>cbfV0K#<cX?0200UK5FX\KbGNAG,1B@[e>g7\NDR4UYM&
Q5X2(G=a)+Gae#Z^,.E6UY,3IVO]6eH;/SCWM^Z6HGCXI.<-HB=C=PSb5ZTf7g+S
LAT1L:^<c-124,VI)_K_))VN>)R.eRcZEU-G]Z(bR<HfEC3g3LASRYf\RU2<I\XM
1.I>Q::NdcIYZFg<+ZQD6@V=,C5=DfKNcBDR&NV&7S=&3,D\0Pe2fI_W\Q;ETa0g
Eb4X?G3N9f6T9-?AJ]&X[8/ffUK(:Y4^.5IX/XV[^^Wb?Pb4&b12Y):=[-OIQA-E
g6cNGGL+SXFd[/M6W9@P@2<=AKb9gU5d0(F&=aZJa^R5/+;W0aJg6F<7Q(3KYDH1
?U9gAGI8A&050FM]ag]@N7O6O.fU_5L^,#7LNF6a_PN_1FCe_<&EcYaVdINL-J4B
072+B(bI0\IPWfPPMXPLa7^4HBNg)^;US#)Y\B)+8O>a6.?VFCXP#]BEHWg?G9\,
VaWWWe,YT=.M.ICT2?=L3IJT/f4&+,0@POV=-L5U@?H3+GHY_HT^OYcCFIMP_JM<
DI?\8@/_+HSF?53P39EA(03#:US87NCdcd8A7VR>,e.->ED^d_90IADR)H@3ba#Q
O@c\gY8BE._;ae?SaAf<6Uc3<67COZ@a;.bJHOaM(?>]DZ0d;FIeOKfN#5CYUNN,
8,H3-C\7S#.9b=/FTU84;>9L^WNAY:O)+PeB@IXCY339P2(TY?J,e_GE_IZGf5bI
9D9ZP77H[7DT>8d&-)OTK-IL<T<9N)/IWCGM/=VF8YYa&gWX[78g]5<S8967;g@L
^Z](b=@8QEKR1;3,eTg7Y#c[OA=RCQ0.e40b+K\M4^7J>@[31;DFdM2K/UNJ6#GB
5@W=O>O]Q34HB[HND#_F\f^/@M,96Rg^A0\3GB3NM&0,[IZa^FZP<VVW/?EV9?#_
.J6;J//6c.X4XT;68QQ4JU?2X/AZb),g63T>-T_96IK^QP9[BFML_A^=T1JE\XJ&
NITH<33>106.V9/QP^:I_Z@\8fV+.gMK;NF?#I)1U_6-R>X69J;Y?S=O,DdUd87f
YR(L99P+]W@S?&Z_QC-GO97]?5TL=,W;6QD=7ebGB5VU9J0OU7BTVL-3M<OL?L]5
@^(-[AX&YD;_B_@E:4?_C+A(+UID:FRdG<?V;aZR9<_NM4FO]YI)Me+AU<;Eg6N/
1+N,d1[.2TI&8]OHD,aeC#Y3=&Nc02-]e1]g\VH#N7=V+b0(UT:X((\#RNRRB89W
a9VW?Ne+I:J=ZZ/HPZVE,:K]8+:1+b,LV-A(G(T;4N,Ic@?:6,>aQ=H4YQKD9&>P
e6/.ZMU3OaSUg99>E4CXF;/JL(TTfF/g.7OR0VAcCLM508+^RJJ&YD/7CLUY?fNb
;+KSV5OC&dfYC[R5YD,eHfQaAc>\cQH=PE5E>:8Y8&E-BY.b1eH7O3))VARW:b5[
<LaO5TV4D0C=aP3c\TPR<[I>97VI,72W]8UgdY#,VN;e94Y6[g(0^g28:HdYZ0I=
b3[V_#E8gS3c;9WV?OefRT)f++^F1[_fffPLJc[Yaa]1/\9W&#<NKRH+?M/^CD&Y
g400VKLg<9VY?#9_)8YfZMGM2K1QH#W+;d9VZ.(UP9ITY6a\YQ/NAWE1cS\e)a[3
af@W7M)C.AW_F^^eMINDAUF/4B,@Z_-cHKWEFGR;7Sb&c;+d,8EG3a+IAK/I7X^B
_-cP^^;4E?97c(T/@807-K>\MBfTa&&N7Wa@Xf62L5;V=^4&[g\#&\f8X]AGf./T
gb)ddL.0[D&@4:29OfU8/0BH/[)#[f1NPcO]TffP0g58b8:0W4I65KVV._^2A[CL
).)S3?YTU]I&MLDeVLVfF7]:E4TSOg81UeS\4#/Cg>T=;X4F#RbW]dJ>M5\,fT5O
bUBY,&6f.XN;AQCZaAXVgVfE4.M?gbJ:7&=>Y)0F8HP4/X^M+NBT5Gg^\N>]K:bL
&-@D.f+YMF7NTF.:ZbW(1)5Y;#5L+>/abQ9STG((aF8E8Y8IVMDNPFT)1Le&M_QW
/M8J3L[1V4->&3b(87XT(Q?;).E373TSAWV\FLBdT@a_;^.gXSb^IdM[M4FCT=^#
+T]64MROFYF?H?)KOaa09JeT.T-\)_<gJ(F,KQO@NQ06GKN2+XO62K]Je(A8V#BA
5Sc9f@&O.XE)V\\gXU;F#>KU[&M2[a7[2PEdFbHKSOM_:AH:#aH[I;O@bM#c=,#L
a?VHT6MXc2g[RL?/=)dV&.S7Od.WG08O2@5K7?5A0A&QHdQVM&g-d?[Ydf)473(U
2,B\Q6WPC,c?+A6>E1#3BJ?0H0e?_[<.BW,CHI\b1SPY(4c^5SZT:<7<JB)]+>BR
KbMNDF&fUE.>c33T)5cgd7:3QAN?ZAX75D(L@=f<>#e/C-5\07-@=CII7DUFT@>I
FW)5=Ka\;^B#5ga=AA?G5HeF76__YZA1FJE=_f8(?CO:X>3LUee&_./H)^\dIY/)
ZL)4N@+LKI6_e)GPUb+BNfXE&057J6PY-9eREO&?aKb-Lg3Z335U6S4)B8PfB5+1
eXV0CW8I?S]>cKOG+ZH;<M3?O/K)_eIV^Q@;AF>3a739;M102K-HYc>6Z0Ff&b\M
LCLD(0#A\R9+MEQg-AI()+?6JV_#\Ad0g]bOQ4M4I./(GQ;K9]262XW0c&4JAI<E
E#_5?_.I.aU&-5^VLS7B0[^3(:7AAT;3((Z+,-75M+S3?7VA\=@L#N-L+D6<VdCC
8X_5:SIN6496&K0#;4@9Ld/V/dWCE8S1J[?=)X\cME(QcK)Z)C:35[1JU/<(FWgG
[Wge+R8,#816,\B;A.N8bE04b2CO5WBRQDd4Td5^I\7e:34Ra2>aFZfLJ+8--:CL
306>PG3HP+QU]TM42c0WF.I>ML>:87:cg1CIabG1JQMR)QO3gP98f;I.;89SR\6F
c?,Je&F&c5[PdSE>5_CQ,FdIb6a&SC-5fUYSX3^\IUdFEcYCV.:>\bGYT[;2e6[H
P_cBdY\?<O)ZO1<b2-,&M=PB:_c8K=0aM=[R(c56+IZK3e4-,&^#C>M1V&>eB0Qc
Y<,ZBAN<D7]eT+30#Z)E-)5R>F\;\QDNc,:gXBDYZKBE0aa7A#[H=K+]#[))3.B&
F1f)dDeK4HYZE&;<I^XOHeJL]<0Bg?X5AHdZYc)C(;]/\X\ZaS>9^.IAa#SNV.P^
P<(0XOX,^[0Y]FV.()^Y.C^-eZ?>WX8WCF0\)<:)H\D_Tb5D/6+HA;0M=)SgO0DT
f2#.M1BffcH6N&0551EcK^XZe=-3MfQ19=83A=#WL\8/ZI>]f?0>@VEG7:e7-9\)
_B5P1gbg/e_M22O)-&JGRD)3D/X]MBE,VST5;8_5@-1F(AAe:aOV];@\&#9XdIYH
[]+IeS1Vc+9fO60CH^0-V,8EJEdRDU1Q=3U9WN>V)1)D030JM\S:7&UL8+A3EP\\
Vg6U&6?.(?AQfM#/KV,C0M>fGa18_bE+BgKf\0I.@aaMB9ZFT_RO5X:F>X\&LaQ:
<_0N:H\G8T,9g\G:^Ie2:MHO)/gWaSI/-1\^LXfA(9AgD9Ad]O;MeYbC<aRZRVGS
IEQT>^>e/@/^-(9;/::&G6?cNHZe=/Cf[\2d+UCL(_B40:]W\6[@U#:cJeP>MZLF
5UgF&PZTF;.-eS\63MBPI^Q2:\a^7d/-)CfQ:,\a5f.H)1<7U=F_Q?0G:H98)-bN
T;aX28g4^J;]MQ_\;B)(N0OL@L>OYF?8&DO##T#Af.\76_8\<.CIS\AXgN-P<9:J
X>>K3[:62;ZRW1V1ISWFfb?I]T2W,fE@>66BZ9OQS+0)d>:SGY1OH(8Z>?aYTYT9
6DJR1YQ&W2bKY0>,d0Ha[0M,^c50>1-:\QX4A[<Q[ZJg@@EL>bP2e[DX(BNaGGfT
&ZUP+VOI\0B_P81[b;2&-R6)C@0NN>/aD0IN+XKOE71928f3H.=3fI.HF]7?=9Ve
82P:RJgJXf-Y9.5Cf\@1V:+beRF9.1#Cg?=S7,Q0-3IRY;Gb_FK3R6TARNc4:=DC
H+g\;I5GdTFUN4N8B-MN7P^#\DA:Y#F]D4-OR&(U>V:,U6?ABHc+O+73+M\dJcgO
K:K-#HKe0@_N)ISE,K&M?RH0B6<cWI5-ZJUX-U[I>Q^#bWKU)AW\gbS,GJ#6I@cK
6<I(E>O9;,\SGW.\66VJRdMI_;b\g1&Uc6YA&-[gIS#-QR6DI>=cKP-#4</(g10+
Sg+f9+[gQQE3<AZ:D3GVO>^9]g+XZXGS&,@]??Q=2D_U7Ua6.Z8O=8OBce1]G/U6
PC@I4NMa)-BCGfS=OBU878TBVY1O:[d/&a9(9QY6X=SHGQC6aVGe._.57\M>1<(]
&B.LeMA-BTG?4g5/F#IQ.G8bOVTe;9_5Ja:RGNFLR.N\eKJ0IN[;[#+F8NVEcg:8
X.(?S))D\DCCP_2,;a(XA-Z+//.^C9^Y\b)AX^<+PKGdEVH1B)c#R6ZVM_HNc;b7
Y\F)Z.CZdVF6=TeN29gE9XbXZJS4E_ba_[>S/U@F34b+F+?f7ENe=CVC7JX?_06Z
6NPe5fIS?gL].(\EGZba<Y^SW\KSH9):;bc@+;b1,_:.[.-gSF[\[)Y30,X:bI?8
6T@&E(GU#32.UD]^(bRf24PgUEfU4EHBW)7&EAb2T[+RJ[WYTL(A,P2V[2]25,5@
#\^ccNY5@]6,>:H;UE&=aCR6ZC>-Bf<QAZ,&B=ENSA1[/cYg2#G(D,M,^=<+<BAO
-P@9dZgcfI7^XDEDdY6WLg2UKF9Y<U0&Q0S9Q<;1F&LE1HWQKVRC70P9#FKfHL@Z
OXPc&gd0^<-c;4#K[KX/6F2(Id47Ke@RX<;Y0\JaOK)6DfM1S839O/PX@8QOg-PO
3J3LNRg4NNPaZcYd]QGQBfXMJF53[e9ICF_&9(9bMU7D-\S5&aA&1VCHVaD6V5Z6
5R+4;aG;(8L3+[,d?/4b.JG0ZH3815)CQM:O&;4&F^V7X^c:=OMS#FSWI)D&A0BU
>FLT=>E&0/)0AMD1N)HHX?;;OE?XS&-3(NN[8=HPK<J4IX^4YDc9_^7[1HZc@ZDD
AZ,5FdQ]S@\AVKWP6P/]Z4;V.C@@9bcH5L.QeOLacJZK?^X6Y>dJ8=^>9adKM@V8
L5Zd2cNV6>03F_cb\LBKg2.M]B3P(GNa8C6\X>9BTJRU0SQ1Y_W9.81]<IF-6Kb=
OFJX2^dGAYbd(\[+:=9XLUS,;11D:P<9VD13QPZ7D:RdgSNg79eY8P-2#IC-T4(>
[3?DYER.53NCg+_bXf7_J)bX<TZ5WK=FH0RF9?E[K__4Z>9.46B@[fU58,].d,LF
(?DTS5[D@D8RPD5FG:C)(4M_J,V_FUe,0K&aQVMdUSI3;TW.7102=gLN:+3J>:=:
9&5M4<d<3[3JOG9fJ&XM-e)@:e_1DTG#:J,)=b4TD:(KZL;5_4.S,]T7UXX^5TQZ
6O@Mf/).9XZJ;A?3YB1[W(fcO3#CFR9ZS3c7T<M8;?1+6D?Y@@\ZXW-?&PfZcCc=
bR0a.2ON(.1OM/P25V;,&c)&f4c:/Q(@ZPe8.^MTSD/?@DFfd#9W.J2KN&=/e6@T
)bO]A.I#:YB<\[b/SY?+5;8/T&W3LZKB4U7cE[27c[]JgF/g-CbKS>.?6-NP=b<P
HZ-M^AYA6f92,-NB5(.Z,GB_B\G7cT9<QMPR2\)HQY3/VVdYS:)5OAdY.a:fJ(,7
ZbeXY#X)KEQ)T?F@5VfC81FeAS</]]\&;TI?0[_+UYe.57PIJTG.0NK/<T::fW<9
>1K6T2R(#CX4/VSc26E<()><(1W12M7J\2MKdWZ+85A:3WH5&K#gXfg?BX(6HS4D
Ve4A/1Z4RFa;[GX@<b=b4?f3Q3Z5:#GL:J6TMLEV^8cbg[+DYV\TgE#P9b,MKV1P
#CVGSTCQD^_A-]A0E_A><C1\e/0\EcFbI5M+EBa^\6IY?;QA=H5I2eZ+)-CF^B0B
A?74fQMK6W5Z1F#I<f&42G/-D-EV;>RDN[:AbH@><]4A_Af,3+D2Q)EKcC,5=6UL
f6[I[C>+g&2b=E-]]X\L<PJ1-KS.5K3@e34&]03CKY1VfW6(&B2=CQ8b>N#fG@PI
^]V7dMDF^6I<Id6Y45>?5(.VWGH4d;_V24V4)g^Oc,]V+^GR=2AB7g^c5)I02.TT
UR5A0Wb-=@TXS[2SK.J;HA]@,KQ/bDWJe&@=@f[TVJ[29V8RbMQ@X.-LaacWYX)b
;XBCT/Z[LJT&f,WTAS_)c.:Qc)]:;<AST\&2V_M(?<PN5^:+G6NcKfTM9eLE7SC#
H.>WFVGL[X^=;V+ZRR5=gWVd1gcfBNLZU)2YdALX7W#a>S8;LTP0&f1,R:GVIKdH
F,IRcU)&Xf\?X;ND8gBE<]2VKaEZGB3_1Gf&-0\=V3e77SUP-b>\.T&L,,.e:.W[
)66cA?ESEQJeg_1_CXL_c37R2D58+&_gT7W_D=V@c/D/V8aR@4Z,^FaAM9D\LgQF
K1gHH?-2#CB\4/:RLEJ-#9.A_-KQDfBT4c,1,^3O\T,BB<D3</3QK(-?gY]^3A_c
+)Y_8c47@&LKTZ6L.^(^fTB)Y3LG7ZJLC[5:JMU?,8gd1f_70</,&F:fN0+5g[LT
IWRb:eSE+:^E0ZHa+#=f]NANZK=d97UP^Fc,K(TOC4_YX3(Tf2-CPgQeM-6H69ZX
Z5P,&)R#78ST@<ZZ@-3.^N07G53&#QIEYbd4e>]Bg<a/9N@\S2LOJLH(GQ9P3Oc0
&Cc3=?;K5RMBe]QL3a[X.^W:7\0e&eS/:d_=./[:dH\&0;Fa..C)Kb9P[8):A4C1
(E=b<Y82\:a.SL)?2^5OecaP>AMeb5-L^_A&UL[cCY<Lc88L;e0EK1gAT)IHL5Z_
?^HHeH7Me63BYVO<f_W#;8eP0A@8[dJ2D:UO(E2gcSc6X#)>M#0QTQ)/&0/>]CWH
bTTVa0_d46@/+[FH+I<GH@-L@QPB5aHHS^HMRSHc,SI)BgaYTS+4-cbDBPUEcR6R
/C3(6KASM+W<G@KE\S_;aKAHYCcR^cSPY:BYW8ELe>a0C1Z3MNK>AWSPI]Ma>a^)
ZI<,@ZTUZeS)M1M_7QSaZZQ?VEQg52GJ^OHQfGQ8)H=.E]g,)HMZ>bC5UL_.O(\5
[)1A5#7L>)B4/;I]F2:-+_K=bWEa3\62JUO:NB.99>.4[]4ZNBYGU,7A^8N&A9O7
SB:C,Ge<aCVPYX0(,]#^]_,WCZMeSZPb<#Af=_MEU7))RMVPSF&1e>[dFdaV7T99
T6E^MW_[XaR99QIF--?\cM<<f<[+PX)Jd7X63gg<SG9:eZNCT_f?b5C,)>?UDgBd
HL#UdbL0N(^fX:RD_#))Jgg9T<:a>Nf](0YfCZ.9R.W[4_45N,bg8([LJ:J9JO[>
(&&XLD>NRK7EQf^g[T:<3JHLS<-T2W0WDS.FBSU8b#>,B?9=H/[<Daa_6PLU0&3U
M8LV<YRZ<^)N?XNd2I)7JAcTI(T3Mb0Z58]Fc[7&6<\S@W#LD0UV).9fMbRK+V?Y
.<<BVUg9HF<UEPS[geDB<1F>5<A+d\3JdJX;L:4WIfR;;=D/8c17KJBR]=I7<N/:
.IIZP3N73CVU;6,>aHFB^JI6+BZ_M&0OFYS/OYH(K_4,bf.>>@Z=]Ya_Q?XO&X+_
aBEH/J6Xa-HQ)>RQM/]V;AN=:JR0OX6)]2811NPMV/4U<9:SA.bc_6:65<0&_Y,K
)@&8[4JZAf>\\CZ<F-(HQOd1P+9&(W21>BD)eO27,eUdNL/e:-&GbQfV#SVM9^(^
\]2@>TJb)g3+\H?GU[dMO\X6+.]d4KA_JQ.8)[^;_Y1MYLF_19.A4)_X,Hb&b3BM
ggER&ARQU6#&d@CX9g_I)5\^5:?C@U2,;L.8^C-fcJSCL86\eHfB+aJHMZ\gd_fQ
W?\>H3-(dNY(BJ^/#B+CGB)/<ZKO-F,RXgA?6L<4]BPA-O&JKb6G;BLa^<^81Og]
6,#JN.?,JCeV>g#W],0e#Q:X8K(Va^a1V:RUSIBIS(\DZE17OHH]dA[EHBf8C]0e
WM>-MWG=6^/UaJ1,/ELFQSC8HL-8&#KF(d\bEYJ22bC;,?9e]N./LI_KCV5a2>AE
0C>A8/[^02c<Y^4J[./;-,G,FJWaU_.5ZVDUc,<O0?J?4[GD\WUQH?GFOOF&(852
7T+5>JN?H;#1TOJ\,ZZ2I=8&:\,1=#5=#>cIQe.\?G7;LbI_I[GD,5AV0)@JICA4
XW5L-WT:>AF8b,\dc)7KT(457eJ7)^LJC^9B?\HdV902;:PO4WL3.\3(b9M/L78g
)]SMH5f3IOSW^Z0gSI5B&I#-c=8#&GC:[&H\X#M344Q\a=#>M[gCBT/.[9?AII91
#&1ZW-+#4D\7<<IYa8BDCGO(,Y.Xc+:<LMO<TCS@T7?gR3\E=Aa9bW9(Geg0H8EO
TPH3d5+fNGT[A,@3QGTK5c2,IdB6I.1PPVLK0HJa=Z#A_(>(R6Y8145G79ET:bFM
@H?K\_?M+6B\8\/,WI;WMY.-Q+X3gaW59/Vaa4FU:5&D+X@.LH<ag_444-W7FgU@
,;f6aTa0aS)U#=;[_fKK->/RQ8eX^fbP::+_+&>f1+D=]<gR,[WK[TGKOO<Cf3bT
aeU&T:L[L.5eA,Ib8P6KE<c\1^,29H.N2([6K.CF12]_EC/0Y,BNCI8@P&/I&&/F
/KJcIce/)CU76WB,W0/d(WW8@Tb4cC]Wc)\7I&P1OV:;L+gS#bTc0^O@;Dc_>ST?
DB7IL^;OY&C=1b9NGQf5?4E(d<#ObS1OW6RJM0)[TQLI<:8QB7#<b9BX#XB/3SPa
6Db.aSf:=Y0)DT6d10E=OQ9(aa>147]>OT\O\DTLVeZ@3&WG6@e/=;WD>c[9?0FW
2K^,MG\15T:_EF#MR:Ya-I_Q_FE-f&>6KTdM9=S<5MY).TBP;M&(HZ2]?1134S)_
J2A.>@,?BARB=K3@=L\-#7M]]H#<]G&4@TH@?H;AY,WLZ,6&SI6BQM;LbP430Z@+
1GK&7_ES?cOXfY9MOD,?5Y\Oa55FW1Z[;6[D_0DF&EKDffd.6\17f@;6^(>#I=a\
IbE&G.XH=4aKQ5<VFS8YKfeCNede7[=L8EAe6(AXE-b/V/HO7N1O+<&gOK2fFW=d
5R?5NCbaUKIUUDZBIR3A@XY.bVcfD^W;1c8Lf?2eC<1ED/#f?f@dP/dI/gb,/5@8
6=^5P>IcJ6:=&,6G,[DUO8a8MQDdFKWRW/If6R53R^U0GZ_[>P=aCQY:O4d=2eBH
C#]IJ+UKfC9:Gd^@DL45-_6^4W7:SZ5KbK8Q7#VCQH@H1d?21EN^#7FIg334a[a9
YHR;LPe-8P20IE[/G);\0C:2[ZSH;;Ub#ULSK=<G.H;C)&[LI-;=L?#>3SP;_,_3
,5:+X7KE7PdVTQ54N[7OC\9ZPe6G#;=\V);;IPR)SEJBfMA@EGAU9Q)-CKQe4]Pf
,g+ZT8XS43Z,\g668/_N+RfC:G]aK1P4>/BMgA:GK46]d;BR?;3H/Y)6&aR4;6AG
6bZ7MP?>(-;Q8^W[J8F>fG/UV\LHgc_=egUcW#3E,S:B30:I7>e<,]b9=8\XYGKY
-EN05BG-9@U3c).)FL<>VP8ZBa+=@98PI,Y):&@W;(f1FU4/7HL&U?4]:@H@:&C8
97UXa2[.2??T_WPcI26/]T9W]XDV\;)6>#&D2;-.71L+a8Hb?O5DOOCB-B>E@ZVe
5,K]DFL)DYaT&KF1Sa4@2-TDX3>H.-SHcNSVC;1TGXMK>UNYP#RFZ#b=I?>TO0_<
I:P>::)gVQ#50IWS,^1E,3d&cDB;^RDG[M8SJ[dXZ,=b>6CH#2.V-8[PH-8I6b0/
)]-OVb+b4T_=bb[C#7f6XUYZMY;)QgD6PeI[;G:g<G&F,5_+J0P>]X&YaaS_,)II
\[;>EA@(^O8#/MRF0b]<CBB+V/J,+A&2edH8XL96Q&BSgIF[WAHH5@_e(Y#TPe=d
E1,@3+5Y3fQK=):Z8^4>VH(KB3J53b,dH1C9+?,LW6RTWR,(ETO3(V\a#c[7eI:0
K@4?[O#-S^>8fVbT(CaO7>U2=;U]M703;R4\EAS,;Q/fZME5QC\^cAS?SFKT\\@@
]_\1H[@a[6[d>_0g13HaHX^8CQ7FT.Rc5\R3c3<MG?c\=Ob5(eKD4,B]@AODYW+S
1;X4dLNdV3-&,+0Rc/F@B3&.O8V1PTdQgWc1[8:V0R]F0SI@d&eETYMXC:TY_66.
-[IU&M6TLI\Pf1ST3_[/3I&3=7#6ae9)MN9La=KdV,T^/QWZ3:S5.;XdE.,VNH/,
-9;ecB&IE_Og,)54GS(P<2U&PBG(.UD@3J9TXW?H/\QI&K1;f(c]BHUK_NaN=SJK
4//VIGbT3R1#V=R1CLTF/2CDMe/;92A6abM(f2.9O&.GML#2O7aU(2NRX0gW3Q95
7V+S=5gYBd_K>f./e8PR9;/9?VA5WU^f/bAOc1F67]^9SBI@fY#UVVQPffFfBd[\
J[KS=LU,YXH2F&@H&cTG1K]DY1,M;@GHRF6f_Sg(9/b?QKC_=9dP[PeO5NO?U:N,
:H:&cDTaBAN&T1ZU__T-7^QN^;aBHO\4.:HK:fQO_8SK_6MXZbGGUeRP996_M7N/
:Z23&W_46N3L9Tc8bd/5&#@(@HDg:KDeHB3e&1R=YW_5(Mg5,R/0A24SDW5Y16cS
?aaHG[2E].M8BRI5Q0_edJ7]a5c7.cO3V9>38^KV/+=J(R?P^,5#=V31-Q5/UQE2
1c9646V290^L3OFUI#a>F6JM^?GIIC(P@QO]-_19c404I_,d-6B.3WLJ>JfFWHO2
]\=ZTZ?-7<-.@f5<MOTB[J@OgO,d_#(17[U+4XVCAf_;&dWE8AI#+FVITZ]YcCdK
JVE(5Lb<IP\fYTLeF/0W@S@a?Z(M:gAe7>V-@_1JPHT618H].IeZLPVKM00U=)^g
QR;UPEFO_=A0a94>W7d4>(=Q&QCBI6-8-<+C?bC@IR+A3VHZ2_TAQb;[]-[DD...
K4(52KY@-,7]/]IfN&HL/@./IILJ_=)C.),G\ZE,&^a#4_FaeWRc4+6<Wa7&558\
;//P(H0@>LYR-GF(eXYX-.FO6^O&TU6CG;/I&_g>dIL8LP[FQ4+/#UL1VADHT)>G
\SCcbgR,(^_fVLRTf.N\-,8+<)>Z[Ie43MU:#7<&Y1\LBecY4:C=S/Mb+.eN=>TN
RD]B\4U4UT^Z.FVUH4CWZ425b[\caZ2H?/6aY30-E\(JA1Vf:gFH#X]ZAT#\TYKB
Ef].@1?P9:_X#^Gf;(5)b+Z-OK2?+ceO&7JY8RN9;,[\;X?>-@Z><,Nf1NUE1?@#
Q?EUU7AL6E1N6]#6/>MZVKH]D/(T16+)c5/b/=)[<QR@;J4?J:MBMY1,B,CI@Hd>
&Nbb3e^OO#.:X/f86dH2R6;Ac6]R?=K&1:c+]:O(QSeN9O2#@FHBdPF#O:_cZA9\
E=X:TPGUO^.+(-GOQOQfA9T^LB^I_86/UWS[OUgKJMgOG^VGI+]..]FA[+bfS54=
5I,_(Z6T(Y@-TJFaX#186bE._MY?eWOf7Na[3^1^Z37;U,^)/IBVQ([c.f:6/#>)
X.I]LZ]gc_0?\UD(+6S6_7X#3^-\4bLRLfA^P(J&ISP4dJ(e,]_E6M6M:f>9TN-0
YD]N#Ba>Ac/3/=+O;XQZRQ3c;VFYeQg]>4ML4+C;:cB4[=C>d49_OE&00:SVLPOM
ZD=0=-X4a#DO,fc_^<.W6JRCg\1)-Cd&Z+4D<e6WB#R5-6d=+K_ETFe@YUeUGFfb
U-,fJV?gXB0eGaW0&XXQ+0BDUFG<\^++-HdL0]9=,:4g2QK<+N?+I,WfB](,&d\1
/<P>2N:V#86R=,ZDA1>PRQMS8V)C0++Z=0D(V&/C_d=g;:UNDE4_fN=G4AJ-=PL[
^834B0DH;D\BWE#JYgHX;_.P6cC9J&W\^\Eg;eF<[U>MOT,;SCK:UU2()F<OQ\dX
GMH/T:OL:&-+G>X</.&9R@A?5de7O=QNZU(@(KPI^0WM0Ta)f3g3#=:2NT/6-@83
@?f,<K4C.]&d7YD[7V+6UMXLN.I3XUCC+Dgf1@<.dL49)9;Je_LB#E3N01(>3:fa
\>=M5HRNOVYJTcTDQ&0>BO(C&94GA-ZVI)>fd0fRDJ&CCFL1+Fe1?1V_0>J^7H6L
G1O@B3-\]1&D_[QCK5.6HB,JSA;_8V,Hd_MJU[cL5XPLA^0cdW)6a#a:aEA^H4O9
BUI:15M+FSXdCLRgaZ7\_;J-?&4EYN\UFe:?(]DM4A=E6QUFU#eYWT,Sg+/cOOK6
SEO^#6gMW1;Z\Zg1KCA_Q7MI]BE;f(abb[0U068L>d<YeM3G<[HG<OB9gWHeDQg-
Rc2d8^PH@5BSbEYW2d2gM&UVI)LIQ[BH1_M\]9Z_Nc1cC^OXY/-6.ZP7\.c@29<5
Y#>MEI13</0J)\.;205+gUQ3[DVNM]__LM2dQAIK<KNfg3_?^IS?:8WbV<K>P064
Oe,WR9I^U(gKY>b@&:^+/B#:bRD-Q1W/66T+]1UAZCe<[.1@/K-L44IR:6L0(,2R
VFTWATH7S]NJ\V#Ca]IYJbXI6[,MaN@d\]M<\:62V1UeDULcOgF;d=7#_,:FIZ]b
N10#)ebFV>?WBI])3Q=,BY0QE/9P8>(c>RRLYQc//A=HFW3N>QW.9/H]R<_PFO+P
-KaP/UC^fQXf0JAa_+@37F62_4YbFe><OY-LO^](P.K)9LUbXFSB^&cY;/fBf6,e
TT?@3Bdc]baAOWZT>A9KgNYYT,eecH+9cGUg8),A[Z&d.cE#[])]ZR(EVC&cWd>g
#0G3&ZC38_.dS,GVeF_dOHRSYWJP-eM><_]NE&7)Ag4M6?(T7LcbP#T.-JZ--8(1
]LfKYUHQ=D.]gMNc0=:8DDF^CQ&VX(V-DX5a0OD9F6MCS6,^XRFER5L>;-e4E-XZ
1;1^U<c:AbG2/PXV4EUcC3acGXGbI<9;.UH.d&7>3OSa=:GDW.DC4A>AF_M1.\Q:
Y,6+dLb9DfI9=L?12)A:N2@,bV[AcGSK?9DA_SO]9^SD?aY6RS<?U@f_dfF/)M&S
?:>5<6Rg&3UR.C<C6W?-Q)D:Q(\I(>VEW,\S(a@YQ(dL^SQJE44QCS_F@FVaSSS1
)1[)M>7c<7#W6J<DWZ1^R1CK81U->2[c.AYScUaTL4LGE1bcU6=aKU5cXUD^S>>V
\/+5JIXeGC5;8@D+b/MbN_Ia_Z0N91W43BF6LJAB\/&gD>eUAaGaO3@b_/fUK@d;
Q2^V.JO>,_8V0Db+>(McNE[X(9-dO,(GYK#a5:ZEEI@L#:=^/&YPK(S2C,R#YccL
0eV<(;T1_L<b5bf_X\L@64=Gg.\_cHc>BWeV/K/P4L&.@f6(gf.gCV\@K)IYC^,8
1]==>163.=;CS7545[Bb4V4#<GMZO/3JbW::#V1Z=gF.OAdC+\+R+W.-TbO(VL(C
>F=25\XBeeTe_GGCNDBG:O?:Q[eP#]cY;;V<ZA1OXX?,]BM;CE)Jfgd\ZOK.b2L/
1M.JK.<>FgJeX.8NJT/O_#T)E7Ea/#<:D[e;]/bMcd5-<#+-.BWaF@L72F825,73
&F0:7Vd-dfS@3VW_bM=5SKR1BN@9QSPRXSaa8W>#E-,&fB/dVdG\]62=f2/QVUEd
MBO:\eDD&^eeUYK94O.>R3@3Q:^FcW8MFUD+DH855;fTE1P+SW63CS4[2DfbXZL^
gUX:=2T.JKCU8CZRT+LKJ:[+WeeO763]8A_a6EZ#2<1&Oa,/]X4D#EC8G:e66O@G
5R-0CSaFW<[B:]\g7+(cI6B>\E/57c;&Sc^KS-e;<5F4D4?N7Mc>KI\]BHK)<X5T
O6/+e(JQ.,f9.deX,IbS9PHIOAS9WFb,SNJd25/DaX_F_@Tb.<a2#Sa<NE@,6X\K
\[/1\LZ,f2\]D[QG&J0SIb6gD&4L],N)K)Q777CA9DP<e:bA26]A)<M[.NNOMTVa
PHE<K7a&@fM]dR,3<Vb-e8,Hc4X/;5UHf#0ESNY&GZ[1X?)EKa<f[@W5G>9R82=/
Ic=+<RaC#M2JGJ2.^?E6d4QFfT;+68=O^(@[(D[;ZRVGAE1Ya\g;D,>4;X7T\GVP
XY\cfM@(-\bQ(>(5ZS(5dY2=<EHd_BR2;.7FJ4[):0aR[N,RW5a,M3\A(?ET?b>g
#LE.=dI-TU((=[)<6dM?LD93/K4^.Q^_9FAH>,V<bGAdP\[@c&@S,<QPYZd.b@[G
V(_c.Y.AY:.^b,I5&B.[CA6J11V1#UK8=3fLcL^&YZ)EC)(C#HRXQ,G7]J+H+36c
OY7d?(IMEDR\^>8FB5VG(F&0YKHNGZQY.CU3d(9/E,)-P#75=,PTd4=E+<G/G1Z=
U3>XF>K@+#:^])X(#W\(g5fHaKDI9ae<Nf(D&#8PD7gYfG]N9K@DL56HAXAFb3;)
1bSWf9HX-HP/Y\&LHeX.W5&dN(#4OgJA?WD<\N+C&>XL8C^.U091[(5XRaQQbN]#
5&43F:+R6cOW?.LM8e4X0D.PGX8Z<-Q8KHO.9Sgc-5GA)X0D.F7#/AYR>K:->dS_
LYDTDMQ-4V;B/76aY@3J6S@LS)A]?4DFI+M;-aB,&IF?5;:]eD8U?.Y8&]8[EK4<
Y([aQDe;[ONHQO<F7.]Fa/7EMI^MWW\K765.5Ye&8<2S#ZC7NCc;,4cU5?B0LW=R
T[\Se1T.W28_]ZJ0F2V>G5N\A7.C=SM&&512WdU;5+U3Q>]IcL4/EXE>)(GGOF#9
0<#P;8&P^)+FcSI.gA5J0\7:)O@,+#eH.G;1?MG.>FVb_eD9Q/8a&_K1;]9T^6;O
ZD=+9K72d<AU+0:TUD2Z_90A+HReOc6\H?[C[F.L7P=Wc>O/5I>?@_)d[ELA5/Oa
]7BGbMUFIW(PdUU)-d3gI97S7RKE9NI:ARB>#78Sg:e9,AaEH/UXab]0bOJ,Zd0]
DVe-3e3e#KbB9,2]_Pg6/<e=aL+eb@=(>6f;GEK]Z5Ab@.F<UDbVS.RUPfdAO(#+
SCW6[1dR,A\<EI3WOZX6>=RJZ:]5^Q<GPe0Ca@LEZU1LVLQ>Z?H<VZXWbBZB>1Mf
V9EGK@?KEJ?>IR^a6C^XOD2#/NJI:BC2E^X&)M@+YeMBV:C)Y(CdfDKT2(;NIQ^a
)OJZ&=?M,Z8E0LC<W6[ZINe^VSH,HT4)4-X2+gLL[bGJYFU+b(PXN6U/0a]X0@3C
Y2cNVM,R4_HTX]PGLO=4#;7N?L[-7=W:SPfR;T6T(_gW4L.K16HB_ESDPgQF5(6X
g>O#@DU^WZ\CL>b8Xc7gVV)-<dGEDdWK5.\0:TDGQbV,C=>6T4@6b1+S)CQAW68Q
.+d]_K&9ffM[aMdY.f3g6K#U^I<cfG[PIIcE\50[83d:Z02PA#LF=NQ)H-\R[YBB
#CM1C];I9+NO/Q.MP79U<Z4DY?346g/c2AGRA=E7<)/)FXO4FcAUGR)&Je+d=:EA
?Q;M6fJDZXXW8;0E[FHFB=.VF?2</HDT].C:J(HSe8gOea<aLc+dL,EKZXdBdM?)
g1JH9<9QD,_B8Ifc8+_O>\HN^afA]42&^,&f[\XM?BME,=J61MJ:[7SKCf58G_LX
/(X,N[cI1c@B@A4249g,3ZMPTIW_DFTeBQY,L>0c:5_3&F^VUd?ZR<LeLWWT?6b&
:OgS[T^+<3YfMZ..8=>#&-2A(^2AL/fJNHe@U9&DYOP;KQQ)@A8\_IY&#8c2VS;:
_eDNXg-7[I1DPV83<B:WS8XG::L(&LF5QdB_#eL6/>V\H,(d=KeDL?1Na=OV8D(b
J6K/TNC]f^D2L=.\XAJ,46G?NWBb#8Z=+?VI>/H4KD)H)Y_+DG4GW&F/7W.<<Z9V
D;&^X_)P\^g7P0Y,1#YcPd]E]G]9bXQF_I[V?_.7T1]MG>3#1+6H35]=S(4=aO7N
&XZe?+GSY#92X;/7^NTNB+XbSHP_OC+E-g;EAeNW3\V^bU#bQV.eW)I/GLD)6I-E
e]HBYPBPLd/25?UP9IcY5PHe,aO93TLVY4a(\a;LULQVOb#GX5M[+g.,OS/g_:_S
\_cFI1?6O(^9c]fG(8+TWZ,/Nd6XXe-+]9T-OD<4-[XTOH?3ba1:RBF>1Qa5Z#P)
0H+&a2ZA00F1(S:.F0S=&;\dG76cCfb7#f323(+S&22)MD4R+>F)E(8VF?U4WU,W
9PJW7:a.VE1V;:+eD9^/>1aD9XJC7F]6ECT0HC#_T(/XMg,^3G6N:\K0AMZU9MMY
gXG)XZ8e,1)f^F/DQD/C]RUXY)O=@:/A;<0A3IAMGR0XeIOU.M5@<50-1(bZ.;K1
<&JeTQ#45c+B>Wb@1;Q@<QF4@,CQNc_6L5K;e<X0J<cAV2PTafU\AHF5FYdI&5IY
@aR\,/G(6<0;U8X@+.M6/&Obb(Y09N#N,d58W:QJG_bH^V7P.T-XX(6TJJVeXS+9
]29WB>NICF(L\#CS/+KgEEC1ATZG5He07:X9;+<-g]4<c+\R,VMC2#@D@87ca<NG
KO(aFeCJ16/>2[T]9)C&PB(cZBBa@2J_PeCWd=TMBK34#]X@1[5M?;_:##+5\3(<
e8BeT0c0@41&U6203))OC>)OPd5YbA1gaI0@E=ZK[&5FBW=N9@X&H]e1\A6.+,-#
;06(9YTP6<>c2Wc9[c+6O6>[XZQ>@=.@#3TO0XR;>&cPNU-4(;SOW1WN1=[G)18+
5/JTU&&(Mb.8_[78>.A]J-c2/K_?XD;H\8_Af#@0GK0-,<#B4]BRS6dd4a8-SOE4
b^?a2?Y81<IBIJ?.d]f,\#abFP\)/:9?FNbS[8K5:HH;#/HC/=Z5^3WeS>[N[<_J
HS5,7O8c,YJ)NTW-:S.dY_5CQ.5D#9Fb6;]Kc)f_\6a-8M[BY#1Pc#RJ?PIBL_55
4G<g0RP859G9b[bSb\=7L^V(<=D,XeO\-<#A_VaaB=dYHM).>bD@2fc.:R,3bfYZ
b-F\2BX.NaZ/#/INY3:4a3TOMX0N/^<9V92-W3a5,YU2ZSN_;_=a1_@+CI/7&OTU
TYJ8;8M>4Eb&KPA_U;]-Z>:J47),Zb;P54D.DUFZ\8>X,c.-W:e&e1SDJ-2;5C(/
6XK:?GSGc]:)BT#CVReAfe]FcQ&JYZAH-M?@83UQe]G1)Jg.=,,/(;\#\#Wf([c.
TFBX;XOBPF3(P8OB.GZE,/WaEe@&1T1B)YY/18Z[;@See<MaDJMb011-bbHI/<O<
R@+cb=SPdL@3gD/&A5(:bWG5+]JB:=#_9@W^IOIXe]]-=g>_S5&-gZ#PB&00a1<X
QcX6,[;//]8A96X7DX;Cc:MHb@Q98N2[<e:dP@+;K#/@Bg#VDVBaBV+^>DTO@(/2
+H[02a7<X6_MATMAFGIC0MD;1DKMS-?6\_)?S(c)Wb:A3H]P1BI_Z@@#fIPgL#ZK
9f;NCIP6Q^AKPMOY^Z/<,0=)gg+1gF6\J?N4IZ9R24/+3bTBT=dN0UB_P:)LHCdQ
+CLRC-AZ=#;TSAA-7D4OKCbFf?#>M5ZJ6b,MdeKJUUa,1ZFDHA0T?X@(0LbbC/0D
>?.@N/PJGH_=Eb&_0:9W:KZ-I@O,D1=_P)7/cV=>WE5VM5A3NeGWFP2A+Pc=7/C&
+JAB8GO(C6+U[]T4DT=W>=14f-#dRVM(36[<^GVX#<A=Ta9RRO]_.c:=a<HPfZ3]
LT>;MeB2>:Y8(ObZXAR:-Zd()6FL>=f0A#_-<WKb5N?]>@cB7AbR;;+/31J^3AVS
Mf5ZMRX-cXFP\9U3<N19KV68=1+TF9<:dYXE\b-(?/&aOORDb6@D1=Y?bQ#3ZXMI
;<49BK>&6Bf]4bNH[feUE^?Rf+RE:)Y:>\T,]CP_9[GJ5fZ7.^c15&FOKH2g>7QD
E9P64AQCa3J8OP9NI#1QC9eWVZf;YFET2[]=&I?121WOLEb;=b^,-&3(3=K/fg;H
TePL(7M7UXRa\U-Q0ee;IaOe#c8#2RGcN@1S\;=PE4/c-VL5).VJ7Z655A)S=T5?
[Z@4UfM6Rb^2b(,ONEHT5.bgU85fAF1QWH#1GH+ZG,VL8c)CK,a,O,]=T\I@L6>a
[OCVX/>P@gZf70_+[J3_YB-JTW-e;#6cKX=)#WAZfX;#0JA\29F=3_LODXf9LLJ9
8)0f:39:+>P-[YIX+-,=EANg?\fSbMF8V?:21WBQcV[G)3H:c,CTO1(dF61/TbA4
(1-_(HI2855VY_5&8VA4I(FCGeU6J_I?/?cE=^D4XZ2P5]T2G.N@UeB=NWFOE[.B
;R84,9(b]g76WM&LCFS&_QT,T2TOYIV0T_]V?6V6(PNO@RUG?N.D\00Z#?XFfLZ-
OC+(2K,S5O[&gM@4IB(W8cb_L;(2Q1>K/W^\@WU>ST:QM8c,Td\IWQb0[HFE@VW0
/;O+=6J7[Z&[S81=\DNG;&XTU(LJ/),Y2RMMe(RU9=g-:E(DZ:.\&2.7\.ZL<=4;
78;Q_.(=V)C2ReLU+\]J3NX>e=6+a=_+TBD&8&gQGAF.-]d+.86Nb-.NJ>Tc26W+
:8ZFH-O/&8g4&(eHc2B4PC0VAG9KdZ1Kfbg:2B3FNZ)aBQ+W^)F]\<NE10KKFG8O
;IR]1V@YUE6CZ.EcLC/UKXIaX+gBb,-.[3,_-)V(_-bV[5(Q5e_Wg4;91U]F>U7H
bY\K^f618QP:=Q?AZX^+^RLH73Z.ODGC+^]VfPO\..@RbFS0Y@AZLTeZa]_&:1-D
WH5V0)cYSOaf-W.+<TAV>8UJZ^=<6B9NI+>SS<-ZMa:0ZA42QE5RM^ac-/:Z?&#V
><5-R12(H1@VYNKD0I6\Y0;0-ga9M4g.7Ed[QF5?dC:76B:3GWY6ST0#M)@PC^A]
G0cBQUf9e++U9\OO6+K-Q#OD)0;W::>XQEb/&Pa6B3P/YEB@g>RUJPF4Y_N5;]4:
684IR2KM#--eSe1B72MAL+\P=DJLP0HP[-aHg[E_c.5(\G/82V++a9#aS;@O#USU
G[aC#FLMID]W<5LH-dQb,_eDT6?eCYF-.1M_9U<_K11U/6/Vb7RcV7)CEU(G7&]d
P7FWd>_A>3//VE3J7aB/YFb33bNKa0FO-QVN.J8a_&1FEP5cQQN7@5[gS01OM]K/
MH[^O[U1S-L?Z-^Z+TSM-KN(2&0>R18^e_?\19Ic&Z<_a8NQ]ZefO&-ZIe6\gV#1
9-_J;7RG17G@[[_47J7LQd/MLW5g[B_A@fEFa-G18?[)9a111fBE=/?b4]U(82<U
fGD07N;fKIgOF+/dH<P:@U+E^fQ0HTQ5)b7AD&97BUfe/2X5A7?\A>=,;b.cc/8I
0,3CP??d\P+J4aTVE4RdRG8;g>e[0,b:9+9]FfH\_2Ye5WUO6eO)]bRcJ?W<-?F8
GG8#;2dEKDI;(DLY3+14RYOCU#e11d(Bf;a+S/f4:R\AE+]F6X,f7U38)E#PA7U,
+1bD),2)4<+^4e-UIB#7#A9@)_7^QeRC17@:SX#[gaZd>Y2R\_:P7S^B0L(EQ:M9
LHO+5&?Jc-^FU_)MWKc[YNB>-d_?^N#X\@-aR,NO6P4Db(GL.BO]]@=)J5<[/RFU
8UB@(CQE=,MY_V9d4;UOX670H9<H@N;bC>\7K3,<_O9&:3AF.J8E=6:OG6_PXKWc
>BA^ASY;4-]/0@C5KOLGX>MEFaS:),TDSXZc2]93X8@C00@GLPH(#)=.[8:K)?3J
CW6_D?eV1A@[L<(1JP\HFHUV1U;]A).)35a@S_D/FZ)6aLXZ+e6@V3\:LUcGd#-^
Wc9UZ[),43D7OHBFa6^@^4H-a7#7+-LTF:00^WK#(I+,1;<c,e;5G3(JN8F;@#+?
WCB;aR3^@2DO)4KU0<HS9N;b=]MOeM/0b40V9K-KMHF.&5AZ7@.OGaJKI2OBN?)Q
Q41_C?IgZKJ3S&N;CEQZB)11XW6L]@;#cf6UF/^.]N5c[[:Z:LC_\-_LHX6XXLT@
6@+)RP[<;E<bZ/RB^g_U4:JH68>4&>JaZA\f,f61/K8N]ZK[2+=LaX)[,^IPODP;
;PBIa.;LU)=/:W.F#,KIJ79I.HDND^7#?g9REH8<11^@J,9/A>>bC4N5WB1a]J,A
QFVL)]<2:KQJ795EXUM4LT<1I;M4>^M,aRBgAQ4?;I3N-D;=3PU)9_Q[eMLUMY,g
Q,<g&J5K6Q<cKJ>470G[O/JNE/1O8P5b^)FdFFce2@1A#\_d:QEEWHVLZd3N/N]-
/T]SZ;Pa+GaURZ1-5.59<EL@PW_]((9C7dZ\N=NDES=57D1H#e;6MEH5G]2Qe2G+
]GP@^B?Y_23Fb\/6Z:Uc[44N68,C5KU=MeM0(]BKTP#Y2_MfMBC>b9-.TI&-N_d/
#MfEL)7)]S0HTfZ8CHZa693<+J[]/+LFPa&\NPGN2O(T.P(GQSHAD+b28HI9c=/E
VVdC7\C@8?NALC;ADc&4;H\/fZKVR#XIMb>?5QXBB,&=5>B:0V/g(7&;I<.<3Cc>
#OKK8;9g>]G8GfOaS#QJ3<)TEZO+FgSN5+#BTL0We7,HYVX>9e=J-([1e@6TOE\4
USf6DdBTT&>Z/59LV=e[57Z3e)U6eVBgYGKL=S/@?IC3?G0<4;XHdM>,+;-R=G&9
g+;LS0<3IF78)ce=\LGCQ_^V426J1]gGIR(a;W7dT[4gSS^.<;,O.CDgYV,cWY0Y
N0+Y#IfdXC4YR#TQ4LgPU^;-#?E-SCb-[X^e.88]:#cJ]Q;GSU@N@I1<HCf<?DSQ
Z-c:VM>7Mb(f9dFcN^_<DSN(1;]#?H;=@BMS#0Yb0]cF6I-:FXd&Yc+3?0f)B0XD
<1c/#Q;f3&.-b-Ne2P)M6LP#8]#CV0f>gP=E83e5T.]3bXJPaXFR9L5^.M>W[5P@
gNNH8PX1S9VU0SK[eC.GYZTbgO)^NX,.JHF+EZb)7a)4>PS.aM<?:Z[gEK?&9abJ
7&Rc/_gP4a8;SJE7H_P[c0@C:cTg5]ZaV[P\KAXIHO8S0g64BaVQL#3(cd1=MAdT
1G;?@,C=8b)5KOVfb<6#6R&(aF9>cc\DBF:=4Ee2N(bI7Rc/[SA9_XU5L;YN:(^D
8f](e3d/H5>-<_#c-&C(SbdZL=5dVXP:L6fR]g1DURR0U0B.FY^,a)@TM\\@[4>N
=D0g#=L0<dWFK)U63_Qg3G6388[_Uf:H^aN(a#T<b98[eP,/beW.U#MX5DDFDU9K
/W4BYQW^@\/PBWeU.=b7/=1[ZTBaLS7cC7aF_BSfR,[E)1#gCQ=[bSS:@OTTS[Ac
0NT@X4Zb1_=_BR8@g9GUZ(B;KcU=gee53E@VI9BJ@C@=VZ,fXH.B>-F6JA1RL\)N
5fGORa&-G#1.7M[15?:C,[;;]:/,RR5SU]GBU6Z^03QNA88O6^d#@=UQIc4P+-2^
Zb-L0b8F(MDZAEdW9_M0gc2#UASAS4B)ffMH8.=<U;eP-fbMG.H5HcX;@O4?8TUf
=e[ePEN+1P5LfgNO(;fB\J5^f6gL._HF5@&##cOK#aL@A91NbK/aYaZN@bXPO;M0
d7#?:Gf+#UZ6eTa+8US&[JM?\;:D?Z/?.9;;O<C(;ZWZCL9++1SK@H<?#6d<&3bT
>LC7+#C=;]HdfS:gA(Z3RQW;JFM1LXEQ0A,M(F9:8>=/a[-G1(YQC4S>Ufc=UHJe
/f^^S+/^-@2D2SL5P0=f<-.b^/4H&JD4a]:?QE\[3A^(fcQV4,1Qgd/.P5Bg170E
/g7W[3a,?=AS.]gR/88:/_I3@UKJED/D/\9gRX1<gb-O4(7-8NCDAM#?gdbZ>edQ
WN2@OB>&2CH.M4\0:U/L?2F,XJTRECa@FIe7[B?D0X>ID0TC>)F?;<_UGK0S^XQU
?@ddT7)]Q7^bBUBg:46_RML+Z4LRL:>9DW4&MEPX-PVJQG]_G@Xae)2A^g1>Fb#/
1^48?JFX1/5gBCS#KM:?6?[1Z,)>T+C)L3X<dJZ,UJS(L_P2?X(&CM[A<+EC\>=?
FUQEC0UU8Ua<GgP@Tf\4VH[0A-SSK[LP5541A(<1>TPfS:UAe9fU6N2H>L8_H<[f
bR#KSO,U#)0P>U)&C_491977<M=8C,0]I616cY]b9FeGEf6EfgR-T)fU2:3Q+DMK
90&007bg.^^HQgG>fKTKQZRU9^N8,VA,/C+F+VVAeMXfU#)#4+?Uc][.^_QSU=DG
4CVPJ9DZ[TD.f4=-OT)>:_-?+c:M<TXQ3W&R8^IG&+^1F7[&dEEMK<RbLVJdESRS
&/F49+97Edd0Bc.)V2I-aRb9L(BKY]gL_[SK3fgg_We<&5:5,SdJb1a6-O)\F/c)
L<?X8I(AVOZeX)Ke6HB:7@QTZ6#_M(b(IESV:AGM4UW@fR/S?7MIdaBXN\:Q6fCb
9CGbIO7>b/Y(e?HLOgY/G(03XBB.C45DD&/A-Y-7b7TMH8EST;\b)RD(UdfRH?CP
NP(@##:&a[1)M,TVGFaCQI_:8B5K/AbYb>^Vg-@#-8[Q]^IfZRd34UQ49;O>M.fV
5+BINVBF=K8F-D;-/c;^257=PVC.6SfS54,#Idd9gQ:;7164-b1LPO[3JG+FVRC.
RS:=OB@HO0H.3ARHR76>LS-K8^HdDUd[aLK69I,b.VU?W0XK_cbLB=e_47Og@0O-
0F,A6+Q-1g7.FYKVQ[:3\Gc\GHAVaSG(eXc6Xf:/3M;&G4+dc+5^_49:-.=(fT&3
=^9-.VGAX3RCbZBd]TJ9&f=a_LXfReaFG]Z6X^Q/B#X5T8)9&@#UC=]dR@ACV:[,
3O=O8[4B[MV#25KEKD-d5e+T/76L99<A3L@R#aLOG>V#M^Y)_K4Pd/8J<EPUgHM4
N5d^g+-VIBV_>0E&6dV=FU7e=>N]:^9d7+)XILXD;Z9SE=#.0.2,gSJ[^#;P(9N(
.Kgc[GFcM:/Q-P/;;V1CRC,bd=AE_NFEgI,#J);ZS9VdH2[Yg^O0I=/F^aI0_aWD
D=FP7b87cFXSHfUS7Fg#L+0((W;V^HRT>6;-?P9Q9K9@L?XSW9YFfTFI430?>\G4
J@BgeV=P\]2Hg+IKB+Z_-KI]d85B-&Ec:#L3PL,f7_KP,e#V+/)UUP5<0P^8>Bd\
U:]6.eIHbR6(&=CddE)2OO-GHIHHF7\U.G+RKTIa8A3WfKTVT<Ta=>5/@\@.,JK3
NWf[RB/bYJe+51K]:8LRMg^G^Qe_LMMD_b,5D/Wbd+GB4dH6F7WD_aP_+R<gd&,X
D^V5MTcbSB)K,==JM1W66Z)-e6La985g4F&HE_HS[=3P-:B4_XO+BFJ;:>72G1-&
;:2eZR7a8E:3ZXgZIGbKf356f49aQB4cXS.D4:X9-G0_/,e,Ed,Z16/\<0[_Xg:.
&f[]_FV(b3X6G4&5R&5R+8RQXK-2.#dX3Pc/\(R,6dL)(T\J?Cf:+R,d\OL_Wbbb
7NGG#-\;2EH0[SY]JfHK]Z/K34^eX(.4VY27A]H(dQbHAYIKRW2)<_UB):>fdF2@
GALTcQ#IXb2XRgg^e9IRLM=K4d7L[;+V2)P]E2261c50.\Q?GCE)gA&YG+FA1N=5
S9NJ6Ve0C,E6T\1Q8(N^9<b-\OHfC5CE/&a,FSO#d_\=AOQa35B:KUgANAT\DA/O
=NAOQ]/(.UU],(G2<:3G-&5X&>bcK\(TA+,<.4C#SE+T#3SbcOY.B].ff)Rg9L(^
\?/OQXF?L;,AA3ZLdd:cIR,:@_MXV2YEfdc&a3ZU3+(2FHZ-)PWD;75T#.BP=550
6(7DPIGa2,>>_Q;SZR@Ya<X&/@7>45Q(T(;<S(E]Q4Dc_B\8X3fDI/<6dC00OL=a
bKX@#KNBT)&QSS=8I#<)6P[<GcM<W^OJUWSUS3&<dRB<3W80_Yd6=06##(L3V\LU
X)5Dg)58cR8]/dHZBZBBK?[=E9;HSdT-.B(U@H20.Q@aJEY0DKc53,-R29Q_/AED
_I_H5@.YU7=<b02@1SfYW,2SNX/=RYK-RYRK:4.F(AMaba2g:H/4^5<86Ha(YZ3f
B1@903W?2JEfH\,]:Ib8UU8Ya<#(.&OFbW?W-gA:[IXY4T5<VgE39f__Y;M9EGHC
8bb<<#A1R1_f9a(1TH7&[[8dW-Ne<fL<0J=?aO,B.DCf=K0G&)YU>4_;&39Ca6[1
5PM560;U9T.N0]Rgg7V1=GCR=YH#?9RBY=#]RV>@0T@1ML(bCJ?,(>MZ;:^-?F:6
,685c7C))\JYXQ_EKdJ5F]/7DFZH9>L,eJ0:H+_2HG2YA>/\@IQgM,N(E3Z-P@<A
:TQ&J0QUZedKU]ea_RO)#T&?,N?]J6P^D>J7H+^OEB4GPV9e0dg<[gY9JO7DCWDa
+0@9>CLEAL7VXCU=+gWBR=DfBcF8f)Y+f7]W/L\8dDBKbYg:+Bc=CD04T<ebg-\b
K^/2KV_L]LgPYA2Qb1W23G&XFHL;46=,Aa<,2XY2K7O7DT\781d7V?N94.L[JJfN
(<>d.(aQEE7R/@+Z5YSE;;>V+]b@[c[[-aO-UIW^JU-HUd[-W8dEe@IQG&E8&acb
S_Hg>/7]J+E:;3G5>WGd[)Y]87b7+3MO#NNW)=^B?;;3fIZ5)RIM2eeUF_B)@b=Z
<d/V,>3Q-?YN0OL-Y?cBbWfgC^=SId3<^Ec#CSAJ0PF^0e\gP/,8<OT2X<VWd5Q6
UPZb]]7QA\.>WcR:AQ:&#WC5E5gb^L9BH7R.QVG:B53UB]3Oa?U7FZ4P](Pb0aX<
.GCV,[>PeNHYTb^?)N[.U\9=PCXC^9KgE:NPH&U1=TFT+IVI?-\H^DYI9)-bU<0I
>JIdFLTOH;S2??F(?9EOZV&+N5J3Ac.8+&I;Xaf#K+YRQ\8;<H[c3>JIET0-,AN1
I2KJ]V4a81X>O^HUHMDYNY9<H-;5D895>H.@/=[@9L8>KM.+/G8U6@&VLSUgCGSB
[-Ea50ET[VJ>4^HJ.:-+gNMR:98]_:7:bO-^V3Wg2#@+efH]bOdS6<&aQI.CUJ#f
?(/CWA^[>S02CI41MB/IQ?X[(GLefL/Gg-9XJZ+CM)W].O@ALg#1B]9?Y?P1\[f)
=S>T0O..S#V10R<P#5#Y#\XZ@-F.4KE/R48<C:Y5Q^Mg7IL>-<WZ>beg;UBR4<UE
I<WT1Ca,GeWHBFfL:82VcD(fJ1;DYMJZ:O2ZB;OgF4[0ZdIU)0XE:?M)c&1-KA7N
3X,bfQ:V<(BF.UH&?,5Q^X399V-d+5Oa]FUAAW#X4Q?0cM)<dM?d8X@7<>aZZ6WB
=W7gNAE3L-JNSU?Jd&a5\;Cb1(>]MgDH=(=FTd3_THYB2Y;>RC0JRMN42Sgf2)VS
?_RaNaUgMDf8f2L2MA=Z/dOKOP/2V3+dT7XbHUN/>/gA23J_=&UU8(VDgQd(Q1fR
[H3g?I_eTdRL(aaTFG0S227?]=A3NR=MgE<=g#\/D2Pf?T@6PZA96[N?>c[5-8.&
RHNMaHe[G^X>YZ?O432X&=;YJ)=[G>D;QBCf&#eXN?]UX@/<7@?Q=cL,/C](\RS(
e9#b?4(0eSN4A(91dLZBgZJ0Q+][W[\14DT6_DcRS0d7B,NG6=aS@.3\cd(1(^R@
I9IZ1g67S1NZcL<+50bdHIWe\Pc:>1cG6_f,)d4:AXROI?Jg(E82TW^+#Rc9<5=T
JY.E,.#VR2ZD5(N6\I+M?/=]@g-bOM)<V,QWC2+2EQ2,DEAFD(V<S,[A61g&0^bH
EOJfKbUX.2[;Q@&S0+5UF&(ZY=TIHK?7#3[gfT_Ug=-L87I,S@8.8,=5f1.Y+06)
(1?(\>,24-QHP-e85e7g\S.d/8QJ;f]bR(I#f<[:<A/>#4N5E4143.T3F80-)Y7R
BCAEbeJ.N8KA46NbO<56c<VdC1VcIU7T93cC;4</=&^d9M4TAKEQdO_K(1b/c^0O
MD[(gB82d/d>/RQb+fW8)9SN+FGQB>B]dKUJcaIQeaWU:^777#.4=KC2<=Q#MH+<
14(JJA9EMA^Y&(D???/GGYW1&QGMV]5:T/dM=A][;\V::(J?f#Y.M&6KE8]/fLP5
(g]\01B:LVAER\H&SJ)bEMB0;#1^JRfb)CSf7CfJ99R.d6ea_([___XXM-4#V@O?
L+3AT^6:Q9[/&Ag<M.e>[+VGgY7B5CTc@d[+,KfT#N,J3\f2B>O?XO>Xf\C79cb/
#)I\ESH@H?M<eN(;>G9>N5ZJKLOS:_<1Q,F\92@@52_aWa]FEA/N).A/AcaS)@fZ
Og(0;dJTU&;POG4e2EKXA2:eQ=-:42^L&cHHO4cP8@DN8gaA.RZYIaT4?LI?.N2C
11)We5&,WdD]CFP?W]_L>Dc8E&QII_>c52A1+&N5BdWKfS=X(NF[;938Xd,e4XZE
A[BO<=O_@g0^B.T4E0)TfX/Z25G1P#T46:;cV4?A-eY1+8COf@HS+bV338JCQ4]G
U63D].QS(a2aT1@1R+ZY(CXT;gHNK+M[U\5GS)[(]C5FCV==&&7Eg\T@<NOdfQCb
V4Ug\)c0Ke1N3@/S>dVKDV?8]A-Re)GJdSLg2ZA0M8O4^^A3SEC^LT(&P]Zd6IIg
GGHBaI3K[Q.Vd+bJ]Q=]I;899P8S/JS4Y80(MBJ_.(C>20)OfS;MKdbAXLD+E7@R
4<NW9(K\GJPFMG0f<JC3EQR#C1XS0KgFNe[XQ0,(bEJ]D;Sb_O)X/af,fC47:G(M
dJ/?UA+1KGH41.4MRJ[A4M#cTY\fT&4GI(<UD7Z+d7<3GL:Cf&O>D\2#8/<dgW9B
Y9gKef,^g<UKFRYL?IE:02B<F;]7MIeL?9KM^ON7E4W1a)]\M)P53H1BRSdW;B?L
P[2<CVcD24XY&X/DX->0(-A][4W4LE>E)#DFc?\6A9(#7#WRS_d0d5AG36ZE(KEJ
O#Q:<1If;1)-T:H&DGHR=WI4U6]+-Q;d]HK[QSAL6fB@DF;dQH30(Jb3e7.36aTO
?7)PWTX/gcT3/G\T:>/^0=>H_BY<L=f]B/GefW9F-E(IASS#dOB@SKBF=P2]/[3T
OVSQ1\^PJ^AN(6M1JDDZ6XO@ZJg?G[IUSf=+=\:G=0=HgEa,_5S@gC==,//0G,7B
e4>Y8.=J)2/5egHW63aJD3A;;9F]>A;F]7f=5NNV4K-6EW</@?Ne7P=T]>2X>aLK
W+b\FIF-P1O[Cdd@^W8^=:)1K+aBGKc5?f2N]Z1QEW-Q]Gc9fI[@BM4RV:a9H&)4
aMR)ABIGHL_/@]dfb.ISfg/QgYK@?bHYb1CQ8E(-^>V#O+409C=c57+/^[?G_W[e
a3SBV30DW+8J-2.U0Z:W><Ag.\@f7J0@M.7)/#V9-.Q>&<SWc&B7L0VX)3O@ABRI
2#-gK6^?B&ZT==Wae?Af<Oa5CNSGQ]G5Za2+^.Y03OH>^IS6_]\e)QD8)ZD8QbXA
W--LO?AD)__)#_8H>?6U-[)3C]8P-Q>cTWBLZGXJ3Xd2Xf#Q5a29#RaaIQ#L:c9R
Y4?ZPP[/8a&6Y+PT@ODC<&LI9eW4,-+eMS3I3F?E^?;ecV/90.(NeGD,g;XCA-6a
X4.-dL/cNI@Y@FT551&9D(+6/S.]g;N1+X@E6RNXB0gWO4S6GYN;Z^@I8).2FJK7
Ga)Xe[EBeB)fV0OSLEOd>0N3_M[8ZLX0Qg-MMSO0ER53?G<YJOO61I61dbb1\96;
UcJS:cNO3g&U0WVa#4fU.-LUd&fX.?&X<PA9P/5_#50H,W3^E9&L4NTJK3+S,6G)
6E^3FM1.-K(gQFd,F=:G?Gd&2KH2IR<W7,b+J?RX?g=]F@9N@-+;gb7EG9b\E<;1
Ba_GOCaJ9@,+(EFLT[Zd4;Nf9b;O;0D0QQ7C&XR2:a[g:dPXI.5#/Z)d.Q494:<Z
DI(dOJ1gMf+UTQV(Z)=Rg&T=b:3Ff0L&F9<=KCSO]<e<:P5g^:?++@=B]HQUG#ET
KS-JL4g#Te/4]EM247H2RC=T#B:#&A6=9Y/89;56Q&<GM=d;#.<H6aHc=Q_CF5M>
2fY[SD<YHT>M:AG,16)<_W=a9b&e0fT7Z^^4:g<>f>W[e>bAMC)QMP81=(<+<8.2
(abA(AG4H6Zd]S74HE&R,&KL=Vf3_DPYV:BR2FaQaP9GG&&bfEReBOS8YS[cbaC:
TX7B9(c+e<H#I4Y7]e4@/4>HM-&_2G4:WWU@e;gBED-)eNLZK,BA94ME)H9,\,K)
LN.TE/OeQU/AZC(XKP+KP[0GK9a6K0XH4@aeM1AW7=PdBfL-7=)R;<[AN+9?bQIS
PFA[1GXAb8cBdC>=E8f4]473gAAYaYg)fAU8f5-X_J>BdT^(LJ]A22>7FEeBA-?V
[H]_b=]]K(3;<H130FA3A:EFJ&cYC6YT>IN]9OGG+B@-_]U<D;AP_)U@MY;9eP^X
<M?2D[-bCP/5e,4ST,_f=[6?&X]_787S5e0cWWfAIYZ9Wdg88PeGUO(VdPW4QF(/
Q&fY?OF(FS]]ID66\MMdB4QMK;<[a?J4=a[F28fJM(\=>a:(\>Fd^)XTNX=gVW7G
F+OEF=G<-<[SS#+[->&#=W0e5R^.V.HB7b5_K:A?9\IGLS)8]L\I19Y_G6.@#8Y/
bH5Q7VbY^5bP;5WV6.C[L(\I3Y/RI#)\JFVHd8ST+UXYH4aT]KHA,aJb&:I\>;5,
)7.0GSX2W8P3c<.FG6>WHgLAQ/R8<N8?e@c7XbJQeZQ?5NS\J7f&da390A(CT(+c
77gF:@NE^0R+&28\@C=F9#c2ZL/J>V]aPZCYdT(:/M=T<5N+4RKD]-6E6BY62?5J
&FBbY9.5BFN9#KN:egGKA_XU=,4;#&W4.Ead#&72C3;P/&PN1FJ@MGJAWUQ=/^#)
)6RV+U4E0(E\TN85\44KKeQ9D]3N0\^>JM8fHH]gTFH=f#BHJ#g4[?dVNSYOfBQ4
AT3+D[KA55HfB2W51?<;12ge&XOaN?9aH.K<&6.VJIXaC6>53+BOC8d8aK>T57SH
]_P7c[J)G]=,P>@2JK4<EQ[.PQ(W)/2;;,\Y&_<@^TDW5SO<@/L^CAJYV,K&=@L<
T^NF]VN#0[UH&egJ;S((#NS)QB20\=,<_+BU_8AO\QLd_-E;K]d1]&Q[=ae1DR6T
+a8A>1JG+J&3c:2\G-?R\Z4M/TeBZ_\9]0^I,/C?,]1=8P-4Lb(O37faX3&@-b#?
WW(MTQ_,M\A@&g>Q2.-?U9Y[.,<>W52eD\(7c+d]g0):W4=;.2Wd8XJ,ML@)HO:4
g_Hd-GP:(TNL3QeW02Jg(8G(cKOW)##9M1H[\:TZ6TR&AG>?aKF-LSD)=:1LKZE_
@M<NX:[aHP94U@MDKO,97;2R,bQR+S,9Z,O5ALO4S6XK5K@fKZdXCY=)E0g#9d-=
U94+5,><P)cUW/XOd2-4GKV5cd]HVVDRM\>[7GBO56.H&1(Y5]8E[4U@V(2[0;E7
<\U\J9gD?[bTLX)_<=HMEX@a9;;7M,#6KU<1<S4fSaR@M_<<6J,DGYUJ.+_N#SN0
M;#C&-MIG?fe661@375+M#06U;e[#N__WcQRTg1L;R;,@ReS_C/a#,,gdNS:S),[
;bAD\WR;K7;Z6QGX3,XaT7/269e@GSQUgQ^NF^a\<\(AYXV+cJ0]d;^Y],/bHYU;
e(HI^@D\f5:AIZdf<SfU#PF,9?:B-b<dTRf_<:^;3#-eA<J9B0BK32G(OFQL+[P[
,Q>O+M\WX;WBFdP+cfRG<f]7#2JG8R#,@aKAb\5I&(>EAWX0a(-L5/&MIL>EgC0Q
D:8C<Ye)TP4.^V3ec8):7HM0c/f6I=cZY8Q3).bVOJgFP@564:9VdZ-gPXRW]bQ4
YZ?\@a7:>1./)N6a+,e-4N+OFa/4AdA=L@Xb#VBcY6G&#NI_TNaZG4UR3BY1_^,b
U?,VWXA4a,Y3G?JIGI8/U=J.3<^0Ma<LA6[bX0CO:Y;Y@<U^g3F99CZNe,1LJR>?
]?H59F^R=5@a8P=BINJG.E,>0YFb@#0_CDCDY.)M+PGdF7P<YSB?R]d6,4bP.QY\
.JA3]WZfNV4X5)+;gID^X;SR7+69CVY2YRALc=fTH/+gSO7?e=(G&Qf1a@4d<&T3
WK#A4da:BXg&(Ne(EAfWO:LbGgTZINe443_?BDFa]6WQ/N9+&UX28H)<;==92O[G
FaDWReQ>U1NJ4DR4Z)A_g\G-g@b=-I&MZa=HeC):PgE2PSF[#2-J&J=&.2-/NFL/
Y5.X[@JW=a1S0@@N6.2L@Pf7OEE_eDg_T=>a3T@D=]^INB0/fZ,d?C]TdFVN/2<0
P@25,a]TQ1>-NfW,Ja\/ARMC[3L\@&geX1C+S<E17@7f>GGJH5:1bNeG7W(:/JMA
;\KU,^];7?;:=Y5WDA3O.[?QRTeWa6O5(FVeXG,2IK?FVA:#M74aV9D=<7>X0c(#
=^Z4>&I\;e>ZAa8d&I[Se]E+7eYN_?P:]=g+-WZ@D]0dF=L,Yf7M;,:+JW<>D?T@
7bGH&#dOQJ21U583bbOWW;UY#@S3=]E2IJ?E+[-4LII_,e\D?@d<_?c#UE2VHU;L
d[+J6FYDYMJ\;4MQ+PU&XOFD_C^=3@Ag\ga#I,3NQ.K+=T\(@gbFWT<KF7K8)RK;
cD@NWE;c<+<da??]CfMQ#UGW&dP1cL[X#?-GLb2<e+O1O)S:],/]IUd;d4LFVWH7
bUW<,18;#8gQXD0\.Q]8c-XbKUQ/9aA])=E-&XHB-bS^YE5EGHb3WY;d93<GIdUS
E(cOY=K\E:YV;FQWLK@N5AA24G?EBc(J(1a:>TNc-.)aZd..dBQN=00YQ^5b^feS
J^D\?GDCWGVR0)aNfJ?P?E=L_d^#G5edMa\I/Ke:Ee;6QM:NdQRYVAI7S^ZSI)-<
NL1/aO(eN&.Wgg.3:Y0Y/3F5C#A<H5OSGCINd<E3PN22/1#,+5M=<+F8Q[@,Z#.#
#,b6IeZM&[(>.?9LCdd6S#[YG7@d5=U6)cH3M20e\g+&a_V4E#<fO._dA,,d83B<
=Y?CVMeM^,?<V(,7ZM1QK.EQVb[8.^YU#Z.97N(GUU[JH-Z)+W)aCUcRc[1e?P7E
d.@6#MR3_._]&;HL:MGBeL2&Ve^bQBYNE\ObLI)5IDS8eJ55U8^Y,G))<(57Q.gJ
g<YN<UG:\-;<1IGdC/?:-U#9R(<08UT70(OHU=V_M_ZLM@Jc@H(XIPZ;eTP8d>H_
G\b3gRZ@E[=FDTd>=]K,5H5VLa873CH.Z/]FY<U=aNP>H36Re>dIGU^O)_(7/9]G
M/LcE.D_=V8-H6K]W_V5R(V^Q=eNK5],g7Lg^??fK:XDG4@=4>TLO]\O.W-S5JN0
J0LOC1[\A0a@>(0X4<K]]ScP\P7Ub#[G&&K9YFPK<H<R?[].d@9XV/VMC(Y4>TX;
KHR/VO8GY:/B+T=LXCL8XV6^_-2Q];<-1Q@KVR-X^SbH<F4:^HK7g?d._RbK(UHQ
&JKfegUS1B_-L7Q\Y50C+0aaN_aV)b@4P0M>dL)//FfZZ[>EB,P9I[(MLYXG[c6;
F9V<FZV(.RTXbKE(ff7IN[0\I4@8-\R#EN8.__Og&B##dJM=VYfEe[FSadM#6E-J
NSFg<3JM[X(SV0P\\I6Qe:e:(^eJ0Ab0Zac.bN\<c1e@_DN&IPa<(4Lc5NCeEb4[
dP+E9a7dbfc\P[5,C1-AD@2gKQ5L05+Hae<=+[]^FKA&dHU0W,adJ@=1FVR&IPBT
3@<NZAJ[)L^D_&L8.;@8cI_16U5G[7Q>V,P<1(0AgO[E2RVJMd32C:d7VZab6(eZ
<QO#bXROdUU[<-NM^J0+d>IOO2ebe?60fTEV.DW+69KdOdK0^PLDD+.Q>AAHGRH@
-_:O=6\#PB((#2=]fY?&M2(Z8gEf@&_Q;R6X8ESZ\RS@J)D@5]cbV->eZcZc)+HS
WRa?_^<DOgRN;]\>ef_7Zd+3-_Q@gD.A6[fU;DdXJU9RTecbdMYG4Ze8I0RgNM+N
g0YF:SAI^O#=MPO=-UYbIL.gI(VUSN^A2IWO-)..a@AQ45&)/P/4&(8e:-?)=)M+
Vg6=V9\\6<77f&R#>W;)EagT&80MOL9@&T/@/G>6M7KCd]O64_&U[7[VUHA\D3_c
+.+K^e,_@\_;_^J<\55&&Wd,I8^P>CA>D2NZ50HJ5E#9T1dK/#+@PWYSU/g?>+>X
D<4RIbfV8,M>)6_f+eHF&QEOHU+M;1K/CYEbVY7fE51g<QIRcQ^K-W^V?]FX>B[9
O&YGVQ/\U2<Z(5D,IXH;__MZ5bGQ?\^F8R-PJ8cdR2^IRL.KJb=L3/eaCQ0@d26d
O2])W\6^DJZ.@=<[3O;.NU=MZQ@Q03d:@_d)IcM?A8[2TNb5)3PF-&Qe)KDOPF=I
G(f<?g5dKE6=Wf.&&LBI.^H4P4WID9Z93?K)<C@dS?/X\0T^g@Tb1SbLR]2SO#B9
KWG.P:^A?6D=Y/-E/Sa6J_TT^@LZOT?81UEVCT6L.gA(P,P7dU/IP.+XQ4P6;.(,
E0F9BN?g:?8D]ggbe=W.>?aWC.eN:1S^<XWd]KW]FW+2>ae#=Z9A-=Y33S7W5cCW
LX>J=S5-WbOg(PX;[+/?c>I7I1aERA2@?VIT^AX#H:ZI#WTN17/@[bX8=cG/M^=V
\ac0+1[(B\0-EYM>P>\@g9@#1/:P>L@g19NVO?V^17N],7ggIYeR#d^3gM^gB;&I
E25CGC7NBEG>2.CF7Y_&Qa+W7L^R-L:S6](=4./eG2D+ZAYcL^Q<>D7eP5gV8M@Z
9?N;MSbKAY/&7cQ7]8,V)(1-VM42-b\YV4Va<2He?J2GQ[4^CX8/_VO\JMXWcgH+
Z^VB8Ob@3)LG9.#/NAJ\AQ;LAN/HL,Hc-((:Ng3a8CN#?7N:N^7FW0QI;HU>673H
/XaBTCD-8(J0RQNABIU?(8KN(Ma]/)WV66V+9ONaf4/c7_I_4V,6K[=Ab6J&dP:]
?#X7Ze)1(d/X=aaS)+1-f81FV#>e,50&ZAW@CcF?-,F5C4:HVD&b<G6=A2g0<B4A
/[=WKW?eAB,Xe@[d6<4I+,XOXaVL1ReAOHbaG6=<+PP609&Jc/Bb(C2e9EW?6QcX
76DgINOL]]U[B6W/T?835DVa,7&3M;FUYB8Nd)T5]I@7X(7L&JT:d6T?7VMJ?25@
&@a3Y_<]OIW0]8O-RJ]+:U1O]QJOaY)G[ABb<4Fa_,A48<,<V(+fXgP[^UHdVAb[
gf7eM44SJ0MIT)&PT@B9<.XNJK<\UIc@A4g-,3<5f[ODZ-+HEHXOIJ1D]+/XMcID
[<T,-Q[4B32FE4^9ea.3:0VM:V+6<,<4;/?gdG@e#ecCcd++-/AIfHXbA)II.[E_
3f>Ie4W<P_^YPL:3FD1M282[0C6;;>GK?^1]dgSLc8&O3?P#BI<FVLZ1KM;K]6,M
/D_Z=AK[\MRfT9HU=1&\Z)DYdO&&WfQ]8#>4;S7],M;D80.&B6&[YYYW_9K2R?Y]
7g_24(19SLTM]:GR/>fP2?_UG4D.<TZ#cFUWecBJAGCP1U#P)EKgZ);ZeA8N,8RZ
9B_6Z+KA^eFgV=.\=UCI)gX/MMfPgT#HcdG767.&<BI_:NKd<R9C7;&K-)2YaC8B
#AGNKHEO-X38WP5.b(6:/Q?\R:K=<8=bBC^XE=Ue;ge?<C//+?.P@.<6)\6O[]A[
,d+F)^[@[G=G;f)&DNe@;2Tfd_8:.cfD-2)X:23+/<eJ/(gMSNZ@gBN0V&>)9/+>
>0R]?.YR;P?JN1,]gJFa/&;T034@OS.V3-d/A,TeA9CUHV3(=?.//Tf5N;^a0NU.
@,B6;;(9Z1b.g3BI>G;Wc4[?(O06-:Te2#??NI6PVY:]R;JVb-J&^]BSE8_ST::P
A#/C#FTf,P]DQ0DM5MVCE5CB]YG]@YY6X4A&;AR\/#S[^,N\a;dOJ9IG/gNdcBUL
de<(W.eg-U#+7+OCY/<[2BGV)-c,b(M2C1BGc/QIG\b,<>0J6W4>.a(c+42<3(8I
XN0O,#fVNHHZ+,ZEcP#64dYH(e-3)0>7E_[Q-[dL(:f+RAeY3\9R8MR=^];I)1M7
<c_]T=T@_^X+B=gHBVOBMd17Z2,8+a:/YT6;ITcX#AK[])a&]^2\Z(Wg3F5e(B93
;Yb)0]PNF<(33,1#O(ZZM27XT-dKbG&^9&,MB;5/gQ6#A;\:?7-ZV[3>/8HF)XUJ
_7SBTd?+TbE47VG4.@Lb&Qb-+6SeQ+f-V\[WQQJOdI-?7eBP/I76^WXG+DU^S/Y)
C90>0P-O;9>2[DJTLa#aBbB1e=eW\g+_W4#=(;T8Y?#F.STMBd8g=gF&(b-Ag^f;
^F5QC2)DW.^XJ:MBY]=^]?:Cb@R_4[;g]d4acQbS/TC1V;gZeYE]\28=7aR,&SC<
H39aRU#T8VL?(0_@P4+>/\KZ\>OFS_V/2fb_T8&#\(K(<TV]H^0S]I:7G..-Vaf)
49)V9#[1[1cU_FJQAVK+-WV20EU\<dR1^HXBf9dF?;U]=:J(-+L.AbOfO8-@5@[^
A6IM9Q/\N2,PEaO/DbS=I3fJ[4&-::Xg:#PETEGBX4F/\9,\HP9?X6-VO-3R^CgG
b>:3AW#\CTe12E1-TK;HH4(WHFIM#Y\VEGWI2,afVWD<F\:Web4>Z_b1_JIXO^d@
Y)+O5(Af>PM9+H+H<cFY&b77Z#HQUgC1SYMW6QZGJ5Ef0Fd:7EZ\V.H1Oa(?SD@d
V>PA?d322Z,=Xe.:^&XPY)=+Q>);GNfVV9N)Ma+[W4,)XL_HXd\#7\OST^c<E_J2
E)I),<;(;L<@G4gMSZ4A)A].g=/MC5(U6[B3=>#&+Lggd]#eM^6S/GD8LBOcQ\?O
F][;]R6-OI_)N1gCTCZeb)S>Rff)Q<eA/CK-@2d]C74ZLDSX6PPMd)e],^;3?Y3B
UXW?]#S9QP=W&5OXbO#;/V<XXSHIL+,J0=M<,=?Y&4@gZI8:X,I.:<-VaMCfe#)d
D851E/Rf3KGbKK9ELQ<EEd7&OLWNS-\Kb.E,GXOOG?4g0eP)8ZBEd+RWA6?J[4\>
5@9R&Q&X):7T=8;c:d8#R[c0@_3H(;<(N+Y[K;U/D3(/[8D[0ZOM-BB:R7Jg(fH2
(KNMQefY;aDMVX?+bA#(GY1+0[[P(+1Z.eJP)99RW&5]3VXNH5]YQTfS4M3>9=L4
3R[=3:fQ;.fZUe8N2B132/KE9gQ40+[4S][)dV30952Ve4+8;2;KgdT;#N-9DC8C
&U=R6Q:Q7NN7]>S?EbLW)664Z?BG[\T2\dHK,\F+D7IOb4+[6U_-71202243MB;#
.aF]JERH4K<.Z9H_I,+(YLCaF:-M@0)Z,G&adSa5HQYDI@A>/TeG^70@286Lc1IW
5>UWC1Y5a=NOPLD+MI9ZI[Q1dR71E\(Q5AS12,#T8@RXTOd>+J_210).@24E&BXa
0,e57QP4?Xf.ZI[Oe=2=cA@88>BG6+X&C8F5eENF&[HY)HF[@O.]Nc.WU>NKC^PA
45=]e6\1>aRB_O7+D5L)S\RFL-]bV3,=M:7@QM8,(>55#+K^TdP0aQR-T>3^J,#T
J#@(_/<>T,e6E7QbG#db_>]B9C?1NM[aV,MHYE:E<1YO9V;?[c;67/\-8aL2#D=7
IIQ:TUg:&A@#g]cbg)B?:eMeKX=?bf3/_^JSNeTB#0-ZHZ^Q?I9VQJ7HFJEVX#6c
(@<.c6YUR#7X&cRR4@3&_15Y]4_]JT4.D/[Q\E4L>@gCX=8.&+M7<H8W5dX]&I2e
/-VADVH2\S1CQEL3dUVS09CC@55FgZ21GHXL,<+D73Jg?)(Td]^dDg7BODVO^@?>
OIHSJ@bgbXV<OH0:KS2.;\-_f6WY0dS++5=+31K]ObYg(Y_Bd+EG]N:+ND=I.\G4
5FFC^0RfAc-I&dc\0Y<:eS6(8_-ZF^GM5HOKT>65dTX?&3C8]aT]N+1.2IZTH2,g
F6=79/GPag24_KOZHWFa,>4>&4@2gf)]5<09;eUG\-&?CI]WcfNg)^dU.BHFCO16
gO@;P3/.4X9YE]+I+:JP3\X?7H8I?(7AZ_K6f=S[&_<D+41:&\/2U0/A+eC680a:
V7<]+.b5B^1?\Tb,7W\6,Zf[L:Y.a8W\JeAc>S@Y,)(B/Xd0MDc1CP?]GJ_Y<MN&
ddGE\c=>[0-KCX.@-?If]GFN?C:F)S^IA2>V(H4:c^WfGFH9GPcb[#S74,?B)F52
[Y[@U6DFFYb3P5B/eO]N:(\;IDR88A&L(TDY__S?_H.<MS,[Wf0R2U.PRXOIF9H-
:+>?N8:>\E<T]YMX6U;-X8<)V+D7)cEUS\0fcLEV1LM2aHF20#?EUS_ceUKbJZ-:
<TX:?dK0CB;.Ug0<<:INQ9#^M_C>[@ae0Wf.>c9c6E\\;]D3&8V4L-JO6OF6\LUF
A8X:C@)=H;ENF9f[H>fB2Z2TN<(;IcYgO#K>O5;+RG(#Cb[2.]e&D,6T5\BFB3NJ
-F?0?#U@3Q9J.]D]HB+V6UIf[>N=L0VRR<?T9QYP0;&e&B-J&(F?I?:_Q1LSN>Da
BCW4:OaBT3aXf-Z\=SgUUbI^MWCg7Ya8E5T1(/C7UK;YAQBP.B[MG[V)4D?JQK(C
G,]H=W2^,EQSb+3:,L41LV/PMe1T)9QeQ4dYH+S5A=AHOJC^c2c][12TLS>a[IaY
_IHQP2VTe/C_KAZ/)_Sf^D0cE,Q3H^Z[[YZHQP9FS<]dTc\Y-T7?]aIdI7Hc1ZDf
b[FL@;Y&H5g8>#ZaK,T84MW8@V8&\DU;(Z>UPV?,ZX.[6<JTe/dZ@+eH5@VP(>dT
feFEK6Y.OJ^&_3]>RIb\<eS#E+5ZDVRH?Z.MPIZaTLLB.P?/a11]3#b?QY#/RRKH
^RQ?-UPA.7\8S^20-[@E+).4]Z/ZT^7&Z2DVc;C4BPFf0,>9OG?BZ@@J9>2H_7b@
JA@-\c^..E2V_X\YXAUcR\,J0M>@:AR3Q\R]d.<S08)V\?@:U8U-6f_/WOJ[</]X
9>ANK&1bWY(f1.b(:;W3ZDa>#,M(fM@ccF?8;[6C_G#HU.Q/<>F.X^(>Z<-;B1F@
=]cF[HT/W4CN_8O;19BE@Ye5@2JcBYa]4a2+5KNI0X<f4TC.=?d)b<NQAf0301XR
),06g-ILWWT3d(Q&fISOO<8J8AG/Y6GN]NC;4fHVNB=J(cW<F^<P1IG2#UEeEJN^
B_>[eYI?#@NFI>V8MEJ2))/3/0[4=N>6F1:WAegPD-5#e07+JRcV6a7<0E(b3BR=
BCJP+<X?;IE.3GB6Z[TO#A03)M^O75.[:-O)N9YOE=:./HUD>^eBf>.b&&gDMI;b
g[c43/X.H;]YX/EN&:[1>K]]ONA2-YT<;_QA?HV;^2BB^IM-Ggf#OZNLG<b#(DbX
6^L64AKQJ<0g/1;4&ORU4]IZXI-,,\aJd2ZBb\\0EJ7V2eLV&HG]B6O6:=CeFN&/
3#(.,b?J?:V[HW=UZfgXQ]Ra63MP4cY;gT9L(KWJI7.15W/;#MRV_=/N-4JNGL72
DEWHL@U8-^B8IJ;=W>#e/M251V0d5.2J+Zb5,@KeRI6fXGY79]^9@=-:C=]S&+;4
4,ZHZ>Z0K.P1.H+Y^dbO-)(=-e?F/LQ^QFMAbFc\R\L0<EK&b9.8-8=HNK((ZVaf
<[TG:-\0683]XV#_6^CDN;.GNab?>\g;Od>M?]QIKGR[bIK&c667a@bABOU^NA2\
7(3:^W]f.-C\FXca)#U:+7Yc#PEWCEZG8>U<3VS)f:fCDMS5OfF?2;Y1bFYKNQXR
b9,ER3c0XWY1FOKB8DeC8fKR,UR_KWZb7Y9WcMUa18&7eRS>E1&<YF8)(+,F)TFF
/24LE6QJ/YM5MT1^0PLAC1GBA-H=ZK5AL-5Ia:DOD#b-2TeE4>23LP4f]R.P]J/+
a\Dg488Pf6[XE1L?7K0,Ae;2KH,fIJRZ5RRF<ZbFLX\4TW/5+7(K_K)Y_KdVE)cM
8-D/\=^=WJ@W9H0>1W>,L/a7JA?f7Hc).gF][29FM^W&ENf(^MP92<(MP7OT:6g[
]ZVYCGA[<-eK;QT+_C+RT-+KNUAI@H3QgFO]QXe9FR^A-EBMZ[8TO^YX6DFL9/1M
eQG>7<)+8U7\&f8O&SE?WIJXX-DBcO0bU-Hd\P\<;c)O,24KX24AP>EM-;ES0fAg
>TB8=(]Hf>P1ba9QU,O&L9><7IV0e#)271@b8e+)XBaA3(8[[+b+Z79&HKF^ID8Z
E)F#U=WH=<UTg8DIbQNX=V_#1Zc\/KD?[QAH/(00)dRfQQL^,\(e#^TP[A9PS0]7
H-5HX^Y<E&cH&>ZX4F^ELaTTP/)C.eLX0]PbEgR7J,_VT#8OdMbWVbd#g>9?=e=N
]BB1NO<M<SIcVV+U9,WD@Wb-0(OQX0]O5JR,2=20@[dBH>>=);:.g+\)2XK;F/Y(
LM16R>eF96=;Eb\b-ZGe[?LXY3+\dF[a7[,V8d\;OASHL5T-)N>>MRB5#=8YLM^0
U/]]V/7AM.f/1OZ_E:E]3S/FM/^/8\JB>BMe<)L_fKBK4[3O+#+PdS:0ZJ..+O7N
YQC6_C;Pb;MHX]YI)a8,Q0CI4Ugb6,HP](49.Z_1Ab@:-BgX1_)fG@\HIPB;f<0&
&7dYS]G;c7ZdF&@=FK:YS7g?EFB.;4VS<OFJ^J7U#MAS?_TM.W1J6e;6a/N7MSKe
R_YNDHQ-3ga];b5DFZRMd&?]_)_[gHba0cG31M#ZV9+#4aL)7:3A)8]d1J_2aE-:
@YcNHcA-DLJ5V139fBB;IXL>a]\/,(/aRX.H)IVW-b=MBH+J1bP?b]<:N@IdU(90
Y+NL.G]<;XMJY\V\a.7+-DUIKaJ+fU9L?AY4)6T^,Uc9+4)[L6=3?/A(HP24PP5G
T?TcC4dC[4(Se)AS[f3L6?]8E-#\(5K-5&e,W]]0CF#30^N<D0)JL5>(J0+O,@_7
_[\cRTSN)-[5JRK#^IUTK0\LJSdC2>&[;32]F#LYDAdgN[51&B::Jc&)(46=(\+c
+,3.;Hb6J1^B^\d,CAB-L;D=d1g6ES[KK\3>\c-.3/X>;a09a/^ad&bMFBg/]7e#
U5&PTOWa?(A&[8Qg>8_/L>a9>]8ZB4Sa.-1/Kd)<]FO=aEN:VVLC)X:7=YG0L+PW
C)/C7D9ZRFHO[Q#bN.g7>Z@]0GUZf@V).H5]7T2V=g@[b,b/:(J+CU)KVAT4Y2+f
Z4KRTROMPI0^He;cWIeLF+g0f^D:bRFFOOg.#.a7.846P&G319LWZJF=/Z_1-KM\
^@)=@7JX;)d+dW,@8W3DRW+^T?S]R&M/);YdZG+FZ,\ET19C.>9e.1FeXKgQb=IF
dae>CTgC#SL]ee:=gd(#4BPb[0BLTV5D8ID?#(\\ffRC,b44bW3,Ea54BQX)OK_.
NH/>E2E0<)@FME^8aU(^57F]]<=<+).C#5?ef.M3Z]RUYHf@\IN;c?5NJ:2W)GDN
FZ0W)dW\.VIfQJIE=)\8cE0THWgP;5Q:]F?:2dJR9CLYNaORMLONP=bTRC@<35&I
@:]04G88P94ZXC]I^U4CMH1-::TWNTSQPU,OZ-:KgQ4GL[;7&>Vf(.;=a?_[[;7F
EV3/2_0J@8+8Y/]+XZ.:KHR+XCS?Ud9/ga/X-45<b)NGeW-M;[:PVGPC>;^-FcTX
R:ERf<IC>OfLR+1-4H?e.^6(?<f;Y?/3M-[N;KF_V+;K-K8>AKE5cKA3/Q^LSe@#
Q^?B7^4ASaXL?HYRee6\c:3GHQ,OdOWDYGP03dN<)K=(>.T&QZEgBaV^FTVF3:Q@
8gSMH-/f(:T].X2(]/Q\NO&Y#A.?&C^@^25fJAbROE:bN<EGfGA^<ZfO644OFNK]
KLXGb:(fO8b+&UJ_Wb0#?R(Y)]TeZ>?>(3EgDWUA]g?BRQcZ;P?Z5>(eI5V)XO0C
a1PNYYGb^&IO_6H&fG)a])O3OMfUV)OKPd78YfA#LQWN>f-2HJQc2-[:?BA,--L[
8^U7+F2NH9C@aJ4-LU)e.-U,5XY]TJO-&\IMCJ4Fb[fTRa>=5JUcSa;IO@&_MX,D
K.WfT4eD-66KMKN5NI)+YR0M_-7INP3K=IMX@,\Ea@4M#FbgHPa@<^dc8L)dB,_2
M&C.9;CR6+RW^LO@3]a]4V+G>P3VEK4BVN&<A7:\(ZWUJ+I5S\SCfP1CON/S>NR8
0b=+@QPOSb_5QN.O0,17ea#[aP+3-FOI)YaGcDB8-=OL0#2(Bgd068OX0-3b=C=4
Z,Q4B?f)CSQWOIYJF4</CaT3JMJ(QdPW9R7YLO)[DRV>I0DCTEO,c.F-9ODMAK7R
,Y&P+J.dMPOFLBe:Re+dI@Gg:@M>R3,H:-HCY?@(K?=47dA2I/<&<f^X_A/d;aPT
A6ARaPd^<.(]SXLZ:3+<[5BYE_IAIK2GUd3AHbX6>4^Y\1\>;0]M89LLT]Ie8.OD
VFWYOFG?[@fAgcG&0<4CY4TXM/42.Z[=;(24b@G#^DXX.()>IZ07MZ(\&#YM11\f
>MW0AA,BTg+UGUP&PXZB:A^S9f[,/S?>^O9/F&eB:Q[gM[4b54?M(;28#SJOf8O>
CYMK0C72C\7Y<(O9@YRV?eI:)HI4-9R&HQT>Z4ePI(\3C;W:+VIZ<)DC/C?M>+]T
^/f)LV7MCRWc6.(?5Dd8PEDO#8[^9aF8[1F/X5;H6=7&H11(NCS0bF,)606[T<aK
LW+cXNJ<gLSHBa)6eNK8[@]L7=SfR.@0V?9>U\P4<UM9bIC0IVdA64^]DbeCB+d2
E.8g&?[F[J)Mgb-+;[LK;:=[3b2;BFbD:7:/K@:7ZW1YS2/C2+0[<HfG]KIHN^>@
+O:f_Y42Y1JG7GHP[+EA.fWFf0YJL#=5KP_=eM62B46Z?cRH]gK3GMb5+PQ0>Lf_
;3aW:6.D+,FbU?1fA\XK,g/P#c+c;BPJgKFSWQ69e/23-RO[FFYc=KbC?TSK(A@^
G\-2SA-AbIDFF::SX@6N\PFK1eVAD1M[c6R_N.CLZ;?/G##,8)XFe)B/aJ3WdF9a
=e+dB1eZ3,YaPBX&KgH/:fGYg^E9RHd#2e(bCcdFGG]=[1^d+C5M035fe-Y?CYT#
(9-=#Sb44_:/g,/+G93GJ]76SGF,>L<+Y/J#],B&;6F&F?@a&W0O<F0<CRFd[:6d
AfMWdK3>c3d&S_?0?MSR(VK338^?^_:(1ANLICET2O+SG3Oa.YY89a1M#6?a<&18
SWV+1Fb>9[^S80DB@@5d@KC2XCAdIa3Gf[>,e1,.BK_BAc^__,4E@)?9WF:.WJG#
J4D;WeO10]H5.I.HFT<(a#aLQ3K,/df71##ec&_.K8beR,7<#=eMFag@PKb@<YE+
I)S>FeRaMO.?(^7CY,_+I]3ee9>5LT7e6,GJ=-BF<N@=Dg-C8Xg^Id&ZF]cF?-^/
C9_]\CO6@U@f&7_A5,@U#?(dSW(H#0N.bC&a0O]R^T;P1MZQ\0?DO#S0#a]fLQ9a
\;8GI<FfS-6=B3=RPTML0?U3E1eY7/G8+#)3L3F=KV:Mff1\V^.?_WEY,Y3LG=>V
?.T.Mg9YIJ=(_#B;#6R.D&ALAVSL.S>7G@+]GWV7LN^-T^;76.LZ>8W)&He])4:]
:0^C8D7a.?D&9=C62Rg^.CJ3W;f60X;[VJbH2S;>6_<ASKD:JXK@)e66AD4Z(#19
6g\QMR^Z:ZR+2)Z,K(HS1Y?1?@1-TeZ<(aF7]6Ff\f4-Z9KCG:b7W,4F()ePXR#(
^X6_\6gF1Y)A(^G#-4OYJWG=N3>7B[eY?)QI9?2Z/OE2C><:]W/Z3]/><J&&[TM\
Z[4E>LU)-FE2Ld/<S7_][7LP_&H\5T9@=A3;#T(?T\MO4^L:6714&]e;ZX.INA0M
ac8aAR104.,R<YW4R<==>cdfER9FA]I:cP5]D;01fU;;8()H8+DF\<TMTcXK#T6:
SKZ<&](8M43K:6._#/RHcMU4O_]GXI,KT&bVQ]4_3&2SV)T4,R.4(b&cN:@3g@S#
^9AAa]U\e8b&?c3cTJR#OHA;&X^9#\-)1gBI_7G3-@Sb7-#\/,:X5g];YJ@IQa<\
VH>dT7)[V_).0AWN+?SL#[V]8-@@cWQ2gP60&\_)_=MY_g7M48;3_KR=a(Y&C6AH
9eE:2?+eHV^NJG#5VC1]G51R1.<:BMfK43GcMdaVBeE8VI6H0:/d;6@8TUbG<&HW
6W0]+7#f++I;+FD]4W5cU8DC02_dHC\9YT,8=4S:I-]1U55:S]F8M4dKLg]RLIEZ
8?JbMD<+9=_@RBP?:-J.b@+-Xg,1cI5+MG],-ZRePB#GZY(?(&J)))OVc)N4<5g@
.S-I=NJL4IM9G3dZ#J2YZ:HXK7\7KVL4(&[9eAV,=T3NKP&VEXd0Q;JV[eS#/U,=
ReX+?cOX(b8-9IN+L98B@7baLa9XI=RXAW+QV/[;1V8Re]-6,.J_^ae?WCgL-[8\
]bW@eb/gJ14ZdGZ\V48bfUb+Q@,[I2015[=8WHHM0G4?TP;AB=9-YET#>GAEJ^g.
^)NDa/WX#ZXEY_Jb=eG55(cB8Tc&1I5U&:#RJ-+ISYd)[1N#A1_=Z898-30]6@Hd
V2WPT.NC3\[b8QA?bF1bc.K)<:eZ1>&b\fQa^0dUb.[]-_<4S][EYW9#<H1[RP=4
5LV(FU-eGD.b:7=L3bJQBb\cR6&5451A\a4YaO\a36dS:@Q54[^8aOQA<A6_I<=A
S8gc-b&Uf9TX,P5A@-e3^&@a7(CC_PQ8E>O#1>7BUTBFBQ5VO4=I2C)7]WU/][:Q
:e\FIOV_.H2:<(a6Q8=L87/QLTZ0^GH?5IfJ:IG?Z8VQYWS:ag2E?N)@S:U6c:e-
,A5gS501G/eG4./54#(F[aeBJ1JM^b/J._fOE6JLA;]7=T<]0]T?NI<#,dS=Uf8b
G+\0bFV9S0bF26I(Ye/5-9(,(&#5[KHCL[Z/+FZ6S[1@57(&VOHe)?M5@?TN[//0
=V(<O2^-M7)J-+/6BE]AA-2eaTZCAU3J#;GN9T\D\-15=W)/Y.^O@OCZYU2KdQPe
.JH]2=?QU8X9&?\fU?=6N\:P_\D\]d7,SKH4X813UL)3^HACP8XYVDY/P\959K&O
8?@]FHZX\/LP1Z,SCC[O,J25?MK]FP-a>U6QB.b/Z,Z5F38AedLU=0V-&gQ4UASO
dY<[OOgZ3.]93OI#bM5=VKHYAccX(_N^CaQ2@G[GcGd(<2NA;6]1La5I1&A#;=@=
LCL[#.:?^\Z7a)>^_^(4OL;RCG<cM/EDL,f^?65<=RJ.TPaDb[GH#MNITEg.DC7.
O(@5\;]6N-O:>?fFBG7\)@/eII6BHWB6LQ(.=894<KCe-?.;+U?bb3XFFQO]WBF>
CedF)U3A;SKE=+e^5/WNAG,^7AQ^=1.&D3LIcag22+CcCH7X(D7>d_/&U\1&0@^[
bbN;V-GJ4<Hf&C:)0L>W]W<O&6N^PZZYd4I00OUbVbGGULN?/+[@4[]/R5HK(CJ-
WTK+71JFK7AOX[D1f29<4=PS-GMg(9QWc:ZH[:K^S-L3+B1Q\Q9GL&\T1cG^VN=N
G:LYKH.g3K1@5:6?TDfNPM3C>0&_B5\WCcg=gLL-_O35Gg3@8)&#B/0EW1+A_)_6
bQ9/FJ9b]V]e)V0TF.>YXe8R@ec=X(d1XH+TU=:A4a(,CF=G4_,QGg>+aG/,1R5d
e-P>d3WXfIQ2-?PP,gA.\R9-4B<^[CZ7FB7X8QE4GH&H->[Z6b6T.(L?g0Q)6Wb-
LU;IJZ+>4H[/E8e#Mf#fZfFf8:8GBH&3Q_0&/c;eUT,PR4)eLKD6)N7R5DBLDaZg
VK-<4_,CBUWXKaWaR-D9DDg>]#;;bL1U.#G1-4JbLRP#g\8dV)D8?:VW-(cU:4Y,
Ra3WU^3fR]<^_(-FNOCSBE#cfN:,XVEX^NTVPP5SUcPeC&6d89;QZ&A?:-L.=5A3
/-2.)fDf\\C32Xgg[]7/TQM/cTV?\a+6L8>:aM08M<C#gB]OWL:@[:2B4#G;LP)&
:1a-^DHKZRO8c.Y+)\Bfa5N9ABdRBNUJ)@B\3PIFcdEF^]>\Q-Z1R]JNg8/76N+c
1NT3c>b9K?N_S7@O8a0W<:FAK4\]NP#?Q8addPFffQFIR4VJ;YJJXH-4e(XR.=d:
Q,:]7S_Y@dAGaNg0QYC03;?bB>4Z#4bK,CVVM[QRCcN>;8NV_0bd<#ZM1?9G6FgV
P;8/F>C^b:MJ6H:6(ZKH)2Wb>IC=/=7R@eLJ9?MU3(D<e@Q_^DP+7&gO]HT0bL8?
>/d[WaW26@f3M#,(dW5#b>AbN?BX2NX9(H_.Z83,2[#[cN^QF)0HTE-FVa8<PQ]Q
S(]=O)L@^14?CW)N6?];3+dF/YVK2,C3&7:FI4DcOfgcJaO2WbfTK<P?7ecM=<?f
#d1K8b9WDJRbI:e)57CbV12CE^EQ[ADZ6WTASC3>^1Wd9OLQTU,)]?6O>fOJ_\N_
F\63abaKR51WVC#M@IQ,TRA@?AfGe9UVSRf<OQ[eM()#S8#UW3M;;=aKeZ[6;^Z]
LKB,].C44A;c2VI@H^SEX-&JdWHGL#I6c7H+e950T4bKc^]_4.G8]_>W3DY/Y2H-
-;56/4\(<->GSNgg:PdMEVb8&AO=Q<_2g>>NH9XSPG>EFaVW]DPaFHeZ+1#TD9_V
++<[<YB1aF3@[-<^NSVO:d/]2>P=6-dW<-fK)<3].]F;XS/I0L9+^@3EB&E[d,\A
+3M:3U,]YC-Ge9IZ[CdG5GC_YP1(UYEUg59@fZEKSS1[0VA^LKY-U)6=H=C^c3c5
f5R93Scd@[,=G4DJ^5#&(TN;:36P-K3T>4E/)#24V7AP1-5R&efKZMXQ9g>:R(>6
3HAXJ+/00B^^aGc]W\)Ac+dR(Gc4V6@FSURXb)<dUKEFM[<UaE^&<<8#KDd7O8W#
WbaF0Ac7&,827)<)R:Zf,5fACg[:6\ZYf?W0028,QGYX,:^0N[116>KOa4:C<LI_
X&NB6;a_CHGcZTOMSe:7-cH+g;\5@]#>\UW0RBW8Cf?^KJ:bKIa?@N(4)I.^[_5>
S-5Oc^L:UFOeV-e0a],_>-Ff^V<P7.5P1Fa0:cAQ=<4_g.IK_ZNKLNbB[/?1@HOX
.WMb(UAGRU^\HRQC+NMFJbF=>QGPJ\gSJC2;U/EVI3-U--JE#M5\,g:\4e13dfM,
ed:Cb-7M=e<#8_;Y(G4MCS/[#?5&>96E?F;IAHa92eBF4(cH=3RR@W_0b8;I\+VI
=EB+M7P@Ld&d;82B>;&9a]TLJ>2_#NfMYd/Vbf9R&ABgbD]NL91Re(SUT8dZbX;Y
&]1;CO/c5[T6(#7FLLXeAbR9AVR3P8>PMDb#f9\<ENNe<\3#gT>Ta9==:CdPK#,A
1>,P(+VX-YPYT,eE3+?E;V+<?13(ETIP<JNT&b_KK6E]X>.3,VQ4W(VdEeHcE-)2
M]bM^OOR/B#+WEO8\d0@L;U]GSOd#fGB4.F<^V:Z-XDe=ME@JV\,(7=e;b+fK]-g
[ZAf1=E-L\d_bOEfC-V@+RD4]II7A;7R1/Q#5]P,52UT61_0/<2[LM;N[d4<HG/U
LKS=72V5DG0^PL6[T7B4@A7(]cC=7X#&[T5FDb[;]125,3/^)+2V(UEY1384ZQQ^
^T4M^<M+>K^_&GHKSVZSJ+g+#NCbV7GJd)&21U,-H(]IEeW/3/[R#TKQ(FF[ATa)
)cN\]d0<UXG_)<Hg5K>4A&SBDZ@YNNg(B]a/_TYTJ1/Z8#Hae/8CV-30QH)/,+LA
\9W3Z])YRBHE?d@Q__EV>gSL@4Ib#:@d/(5TIGb2gW55V#G6TDB^W@-AZ0]a1U)_
]B3-)TQ.C@c4W#aA[<EEEB7IO\/2X@eaG)WQBe(U]B<8a?>[CRH[OD)Y&:d:>DEZ
JdD7D#2O2:[gH6Z^#Ub0]e;DW-VUNH(?:M):A@^d\fE)]^T^YC@NP5PFYaJEFWe/
B5EB6KKdTKSV3YZ1J/QF2_>MED6W8:#5Q-->\>45-\BaB;PU;A7U(BZ)PeBG#5EU
cIGea_P@,STcXRSP1O9<4K+,4P8_)gTU)a)Y&W2c]gPDO013/BJgXRAE<50ILWTe
Z=I2)<;Qd=5W07\Z27&K,^,-ZbX2<72M1dZX^O5YB,^2dcQM>,I,N>,[VVUc;Xa\
0[+[FWZ-V1_5K>H2CSZB:2Y0]RL<,4OO9TP5E\M5;LFD8b_]4W:9Vb.;OH#G.ec3
0Y:JHcA++]7Lg9]61CDICe\d_#gQV@d+P[?X4^(FG2ZD=L?@C(f3#V]fH?Zd<eVV
U.+=f2O(f98Gg;R).dc(A):;gAH13<Le7@^&.EJ>A\eI@U/O#gCNO5&^H.Y;dW]I
]dI_95=5LYKAJbNE#aeGcdL/8;P[=Y)gUD_M=R=55P5X4:[NV(O6@I-;X9NES<=.
e?</AD4.LcPH7;SDH<+1#51X:735a+9CCODH/2S=[=N+ceLW\aB8,HD0PIS=JR8V
g)YT_URQJ18<-8>4g03Y^)QKCaE+4SA4NZeE4X=7=3<:XX,?af2df].U5P-<15[V
5&W2(69]AH?#:I39J\ZcPQCa_X7a151>1H>FX&efVWP+Ke57R]YQ=TDWOKP55^Ad
,UZEDgSQcG\eNZ4gWe/cV?f/VV05/B>;2O:?)8:VCO7N/d^M.fR4&7E>Q64[(WT[
]X.N(9+EAG[bM\KWFJ:99GQe6YA1VW\a<>R:H33TR8bGL^=Q/X\aA;F:a2))=;Ie
?]:B.7&\<BH[?1,bD@@:94Se6:K8N-HB.._6;6X^A.K9PZ6c5R-OC:\[AXU_?6UR
?7.1I,XG4/6Fg4deV?:2K/(OJ7>Z^TF3beaA@2);TUW2Lgc;:7MQYR94FUVKM1d(
_#J1B#G^F_M=X0aEHDQbB0(H+:GXUb_.B3e@cXZ3Ne9>SMAG4CABC8[L0069O[NL
=(8?4?3QTF4U;,>T]de^(HVf\T\39SQB8TSZF/D<1EgD\:8FIY&F6R:V-\Q3HPMU
+ADL);U?4fgdTT/6#Mb;1.^>S8EOEGOVPWSK\(/_07Tef;]Q+f9,F<4_fHSU@,9X
d^N4T[YVg>GXTAa>#I&QL[HOD[I;/9.V<1,Y<B<MHJ2:@[Q/F62IN1f^3;_PC[\^
N[0K(f.]B(@]25<Of,NSZUX,D-;;/F@PCHAX-->98XbIRXEO)>&PLP4O17<E8&[X
3E7dAW]aYccDSH;_a.V,0#@&CTO74HD-5f,W\[U2J^JDL??bTfPK,QbWF:.(:Ng0
<c2cWD#-&/PfL2c9?A\^6ENfVb845C3ebN1d1D#+gP^P=H9K+K1DB@QR+(a]Ce:Z
&S4Z)41&HJOA0XN#JB/8A\:6>KQ4CN6\^2X]a6G0G\KBc9#8L0AY;\]S95<F3R?d
V#d/&,8]:dQ?fX3?b^?>U_GbOV+H0ZO8=GaWd\^7&8a,RU,d3\+FbEYFH6:cWf)(
P@Fb+^OT84,aNIGDOaLFW4.J;9JJY;e=+<L09T2<6K5bVD6gP(9]RG),0^1ZPC(,
A,,+VFCILKTR<c\;:gPF3-/+((5ZPNVa2->LHHRe?GZ5@f[e[LP^cfc]CcSF4Bd[
7NGUE4_)XU#H\#5=IgPf\CPDX@K#J6f2US:;USeTX+F_6;30eY?^/.Y8a4H1O2CG
.JQ<,JD#Y)C>]4e3/aDSLUA6-cEKDcaJXfI=/Vf-WZ3^G02+Z0WL>G7BKYD^[HLd
B1X^,e8^LIaHa//Wd?C4?A;I[RgFV1OUC^N6\/HfZb0SVNJ[K:N=F6KAQULcZe:F
&WQg<7CE@3N=T[296<(OX-P-DD1MY=Z,Xb#@6SJ1>7\;55-CCb-GP:A]1?R&3WBC
fK/>R9##:+7<J#KS:DMfRB,M0\DU#QJG5-),P;,c4E/8+-Y)AP1L6aO[\)1g=\VC
L+Y<NP[RY/,YEYPZ-CQ.9M@)^WZ9JO-/Z^P&:g(a-bX<b(+6&,A5FI^S4?R,7Q>L
V5f46P.N_L.[a2-Q/6TcB?4CZ\,+BY;#XbXIBENND-O,L[5(>F12+L8@BC=K8(Z3
A<L-Xf^W-TLT+S.c;[KSBWOA:LS-Y9O3H2N6Df?]#<cC<Z95YLA6=#.\,EE6I/aa
g#LZ[3?&?UVDc&XKFfg^c(SfgEI#PJ,L4=QJFegB??.ag#HN(O4QQ6?YH;3[OHdS
SP5UF-2;8(9+,1+DY6W1R3WWYGI.:WA./Gga<[1U;CfgH1CVN8b68c]UJg7@&JD/
I/0-AWYd5+W9+JV=/fPS:2BDJ&b^Zc4c@2g.W3,BLWeW9+Cd-V.,2:[fS.\XdQ@/
A;G(2++;X,+.8cfPeOAG[]^X@2DS?9D)#d599dH;f@LaRX>@(GgaJagQ(,^:[c_,
g9=c?#G577Kc5P67PDLT/[T1]C>C:XgPX#S8a.V2<LJ3LZTe:3cL3TXWgG?#;2WR
Hg#WC6(2gQLZ=/:6X4I(M/\O]=Ie[\#3C_&+UUT1[KKA/SXVP3CV5/HH84NaP.I#
]QKM<G2P3>e3TGYI+1_4g58_/:23<&0+,\?[.Cf=F1@HOU=aE(9HPcT@CUb1ML<3
6ga,Ng&94#:)59CW=7M8\8b@2[6NO9H6=KOgY<J3XeHO#9YZ9SIdaNQeGcJ8fM+#
J9e2_006S8+&6H]ae+OYZ7,aUDNa7\\U2a^87W(H0b9\/#EC?F0-BKU-6JXHH7#5
U53(VgKgM;Je2?=)-f,<?I2]./\R@3#41_S#c6D3H@(Y;6aC^S+7F.TdRE8]fOW5
YB1@KSVfWRELfKM)-0R[SD<?1fNDS1\0BX)/&?E_gc)YDKQG(U@KM\J(W/<(@(4(
+)?4SAWdQLN=g77d?V2?c)&cYIDZZ4:KNCVdKGe_2#XTe@9&#\2E5=1b^IE:R98c
5VHSHQC=J^[-YGAX<-T(.^A,<S::XQ8S_B/\4U(Z]6<6AVOSWVaD,B9&SREbRV,=
5]_X.&9R\+MM/:Xb(TK9V>g[Q>?4WTAM=VEAQ_W\HZM<;d.cR4+9=A(8/KJE-C2V
aQ0]7b6B1KS]IZJSH28=6=8ceL#T<97[7gTW8QbGI_T;[^:7HP8d>P>;dWM6,K&J
4Y5]>D8]ag#)T^aFZ,DIF.:J6JZ7S91IC\-CLgY;<E3-M9#AVCA-3GO0]^BPDNd8
Z,8(Jc\Qbd]D&CM)Rc2,;,BGbVJBH:bB&E2VLW?KBSAAZD^#KG34-L6e;AB<:<T(
7?<P=NMcXM82R967U5]FB(S-f/NM>@7O/I\EL;N<3c[eG.WLW,&+e+G0F_8AJ4FH
_]3YB&gMVW,_S(PB3;;H&5CTagX@-=gKbX>]CWYO<L:_bFR)f3b7bK)PQgH<\_25
D@]afYYNKXQXH304O@M5X_N.Nf>/-f2^8+SGRY=87L7^,Z+5aQ;O<Y=M.+-1]:f3
aXY5KD6Q267PRF-NU0faMAE&LN_KPeTQ,LYGa]OE8Q5OO2#IOAWMJ]LJ5:?dGQME
DB9g)D:ILVSD8B4\]L5<I_^[B=/DL6D0XbY4-D=#.N(_;9I<J.e]+8WSDf,I;D=K
=Q:PZTP&A.>2Z?HR4Z7fJSeE34&AVY8D@O>Mc>Y&^:O_/g>K=e<EQ3-aS+9T,OQI
]J2T8P@3GYBe#C\#^7@(;eE4aJ=C4YRN6TD3E18S<ggB]PfV[^cHI=N50c+19;8^
e^Z\<-LOYD@&<&CE<<M<bcB(N01I7aVZC&S-T0UJO-I5cb-CU4G@Eb@4BcR,J8b3
^?\-1g2;:;V+c3dP[gC,0.:^4P(+&T8f\5_TKP&/6C6YGb.g)<d;AN)?6\V(IDb4
^23Rb96QM&ATULI=(ZN3X;Bf-MMAEI@P)F8#1P7A,?RF8ca1:P\(SE,,]d:-9QOg
e8.J4]^+X-_LT+5Hb]\O;.M#_=87HR/&=_3f9RHB^:IF/YJ\B03@2=b8@I=_DKHL
ST6QcSb3>?.g#/P4fNQ=;\WU\a^O>]T/.[3#S8J1J+b\Z/QW#c95c6AC>e?JSRa3
IYXQAK8f]Y[E-gN-bf7\M7dCO1THQ@ZI+c4\5cbTd(@^H]@4cSS.T0=7(M1I(=UR
E7B<1LK.7#?^8_:3Q_V21EAM7V>S<+cbMTMI=1SB.,3&>E924.f2;J/bO\94(LWR
EV92\).NTHW9J>dd(5?;3gM8Z4X\T:M,P1;^H0HR<BXH5H[e<3-g^CV>5/<K0NJZ
RCQ(H[&L8[(@MO:>-UX68<OZ9KA3b\NGAg?J+?V)V#R>322g,>/RabL[:LP3K?5N
KO)V13>9.#264&-B9AT_MPC\AM;I,fDPb=8TMLdg;+d23_DCB=Me1R18=]\918\C
T=\>NQ3;+K0@V(S;@U1CQ=)[J#BPQ.&+ZdZ\SaBfCL_46L;TFR4eWfPK))8\1&>:
M#R0)6dEOWHA:Q,g-\cM>0=?VLK,U2M4<Bf+:+ccWB2P?5eZd.XC9;DA&.K@LECD
2V[DW4_IGH)ScZ=J__-\cN_C0>SEf]d1;\\1bc6T-,?6OI[<K7F5;KPSEa6YF=L7
P1Tg;54XP-ITALdQL4;Z27_=T7:QC0[16FgRQ3LI>Y]BZ7dFTIMW?Y-Z?W(b4F3/
ZVNU3L3d^-f7IPd?\ZB95XK<d52TD#f.AF.A01.TAc>Ta4-V)XT6@XBbKgNa)T07
-SMK;&cX/N-=gP]X5d[dHLSC^QTK/SH7.<:6_[:9W&gPZXB5\:e+U4LEP]0C.,;&
9H,;0,Q((Q-BK2P;=X37Bg/Q,(,.[FRad1Z4C@.GK^##+4G,HPe:9P#ce5@YS)bJ
F24\S6dZ-&,C2/RX=b&)E.R_=Gcd@I64(Z_[?M+MeJFWQT)egQOcA>c#U^((9+Nd
gOX2\J4MPaG7Za3(H9;@eBU9/_C(DY>Hf9WC@;;f5bUSB\47U2KQD3(?#CEKcTBA
J/W6@T6WBO=[&2BD2IcDOP)bfZgKOPe>MSI9>?Hgc>.7.F/QMaG9@^Pd5eAX;e40
),cU6U0[<4eCQCM1G=_0,a=[G&@W[eM&NKE=67g8?:=bF/7>W[3B]Z:bT2e0aPPf
81/V:.L5J+#?,H)aXT5B.W@L^J\G0>SPP[Z]YGOE1^[_S=a]\XgaXE&(XebD/J=N
IT[&CZ0Y^:[.UL67T)(Bc\),#8\/K-X;:gE5C6bL(TIS?QHcB_AcBY/F+]]:5KUI
,_7fFN>,2e@O76+0:6^56[Sc1XRcC:fd4-/0?G1B-C,[4VHG=eTQINb1;B#K.=3W
K5K?#/9AcV(_-5e^EHTTedXdXA@L#P1>[IZMeUGJg:(FU7cJ8Rg3M7WJK]1;0W/Q
>COOOH2,T)gZgDR=#fJW[#5Q=<e[I=)TX9bNKc87[MQK27E\)DAO]L&LdZCDZ+7Y
XNAAW6=/Y14C\O;9O()V_&R3,ID#=?52G=+=CL+9KIXcV05T0@RO9OH(W(g;PcXQ
RVKJc_7IZ9#FB^[f#QB2H9/>69@fg9<PT<;+b?39Sg+-JR]75B9>\P+FgA,;L?>T
D4aIBXZ-(,E[>-8_bAS_>KT[Y_@2CE.:,&@F_aDU;9#],GaV#2eaWI#&V[7-E?)X
&D<ASK@O2TJDZGY2/U.eeS]:)550;\J..c1<[]Ge/Z7Xa4J)Ue,eCEMO,5BU687B
6dD@5@SSC(c2?U3X/-R>3ZYXNW0OWX(B>YE^;4XZXcCc,D@@^fVcfAPaa_Gb[#XF
@>+Y\K:RP#H9R9LL^_W.eK#OW[<:7E06?LIDTOL2=Y_2>eYb#X+<1U(-<edHQPP2
dg\K^5;6:,ILgKF;e(RbGTDUP-D-_.c_,3?1E&W_>].^W/=e<G8M9fC#T2/22JOg
R2gWY>K]?,GXH?O;YWA/)-)d0TRX+VTc\[_A5H1R<79WfZ&ebVEE8-&QcNa)UgTR
L>[Q3R\8Z_eV4+@C6.UF4Na6b,+V<24P6P^&7_a/YcUE<Kd-CZc69#HcXa.L80He
Y8H#c#DfK[2R6gdI4)>&MPe/#4PbeRf-C_;R4>Y/\bOe]9#QDD/3RLH_YXcVCH,X
f:;G4AQUYR4dQJ2YHN8^cZgFT/#&5FV@._-.FGP3bI-+Z@LC-9Q>1=P?Q5PH7fH+
cb(C[7E/fgX1ZeK3?+L8gA-GZTeJ.>&#a8XDXdc1_eW@O,@ES76R.T^M7X49U2.-
ZF[L3+O_6(QXH_8JC4N63;GKGWAb>9^R[6Rb0c&7Y#>;3,4]_EfN]LM,d1Y471?@
)JBaA;]U;VF1V1+],E^17]gOW_9DMeQ7GL[^gTW+PI]V&6,]YgW?)&:8F(E^D=:d
<Ae7?J7WV1+CL;4-\\W\e:QPSa8QB;Y@O2Ybg8W6bTVY?NYcQO^=-=3&K-RS\&.g
FL\=:dFBCZ88>H^S9)FC/f2JV77<]@,N<eM7J@.8C7\#c=7eeORS9#EA+1X3,;91
V[[GYKR[bOg-?#P@1Z_H+=XHC1XZS?:ff4X?6Y=,C(#Og1P9,Y2>3P4/;D-2)b3T
REX+BT4g7\LaQW@AD+FS#dg2_TE0SHV2D/H_+8WJ0.+91JA.OfRHT+/QD(C0fX+P
-A8]:XE:-;7TIZ>^\\eUe:,\689K.4aXO_3Q[9AM\]3=(=R4-\Z9cQf?5/O-F:#&
0\7JY?:.Q76+^^.cdc.#[&7K=3VDK+Jg>O/MI5H/XAX_[@=Yc;YMdee^/^-gd]F?
WFP21@)O>V,c3UHH>J2bR9f,VHB2Q_)K&_G=e-f<F4(c_7VJVd_JZf4>P3P(N.0Z
GZ3:^_bfJe704I4(XW:7\KVPCX:CCK>7F7a<84/_CbZ#eUJ.Y:_9>71?5QTNH(3/
/UX]b)VL@Ug^SZYGRAV9.be37ENW=YW+be:KU0)HP3LW.5N>HY=)=OCNV.0:G<RV
THHI3H1Pc^9d?GDgO7-Z_L(SP11N>=D/R1YW:-6Xa^Q:d/:M<(:1b;)Pca2-eW)[
KaTO@TQEL)M(1)U@Z2d3;,5HdcL<TeC+I8;);JGZZfB_#TKe^=B-#GP+KFF5V1Pf
BYJ2L03TLgA>2Q;.;a/#]gePd@^@,eBR]4:XLP5\<@@)Q>LC_3.U<YV,dd,4FI&R
?U]/#R)c[^+K),;(=-,2Td2)PGdB[f8bZ=T]0NE0X8T--JW&IdI6R_I^bOT?f75/
aa>.9OVY/dH>?HAM/53L<8YcT/XBE6OX4Rf2/Y[g.@MK0.G9f+UH<f].JWaYHgU4
).fT1EIFC,[6T8YNOT43N&N.&H^O^4&0C3(XV:J,<5?,98PaQ@3/=SK.U+KMOFO[
9J\0-BZV8fZLEJHXE2>\Ud)=H6H2,O[,\IAF=fN:a/f6=,I23cb4Wbf7?#?RPP7/
.Sc2=7bCN5([TI/YE5?D=(+LJ.7.ET)gV7&E.\/LZCW^JI2M^#&L[g;^2:;GcHd:
;KFODKU\Z9]0@XGX5DD9\2):&]3YLV4(D?)^.EKc#0dH3;^/b2]FBUD>H]dVD#Y&
N5C2AZ?,57I1QLQbZdFZIV]+0_@:cIfD#79QP;B((/B#9FD3Ha2-0D^5R_E.C\^G
BF=c,0#YT:UcJWL07C6_GB[U4R[HF=E)-6-LGBEE0;7Lf1d>I=V&D/,IX_]/2D[A
K^O+g^/=gXf8U@GNf^-DM+-1=Z&SFX;,e7HTB39bW,G7+dWCL,9JbFQPdeRT+8M:
(DIKAN3U]:]Q1YQUCR.ZB_.-MdFLg+&gc5:=0dccE0Sb9XF:;^dbA?U@XS68DONa
aA\@8N6J)TD]C;L?Pe@8.=VBNR^\NHLg,g/6?+WRJ,SI-MMWV[CI(Q[]F/&Xc=dd
GL)ZE>RACOb[9>?OH9FaQ;a+6GObgD_+d(MH<cgdZ--,PO8[-0.M4[3+Q57aJB.3
<P9,@],\>_)ISQ=[N\V:Ee<)NQ(d+Fa/J#9W>eTe0FIg9)0W0BHQ<0J[/KL9MQ^)
g3deg.H3H7)Kc>R7FZTNB]/QIBG_c8Y3=WNdNI@d4g>URWg(9WMH&HPa?_RCOF?B
8ee/?;;O&Ma;2=d:;G_4H[M-6&[eUNA([K@Y2HB4T7eV]X8b7I5,;Q3_K>3L^MX;
U^\N:>fK8S2K-FLKcG\:V.B_.;+&,?gL>TH=b:3>L-+.5&?CCSg,a+7O@65K8SM6
9(SgPW6\Q2aC=?D-:QU0#aGbFEH8f73d31AMQ/KM.G\BHe2LVFEgPOTcIaVbJQRY
0\Lg_/]:/>X?eSCC]7>L0;:,CE^\E3ab2g@H#4<H8QVMU-@C&L2G35O90dMHV7c9
EGA=g.d8Y0J/Q)b/fE@3SFeZRNdGII&^4)#aW\OJ=LDMM2f-V)]a>H;O:>F;c#2]
3<]f=1fJK+@[HL[=>2[>+7VA-BgEE_?KZ.d;a^cBE4MIJ&bB^(^8/^/F9/,/]XC^
ab<A1DQA770]0[e[FMeW<#a(]8:2fcWDX<7BaKZGL;EB(S>-;L1]+1R/@Y<G,VcN
]@=RM;W>c)Y)_5L_afg_XP=IXd\IPXM+1;I[RcISI-PUV@&a,gT6_a.Yc-EJZA6W
8+@,eTI.35C3.+aSgff4Z\_.?E_[<8MK5KgL:ZZIR9V)B;3dLY]L<a/ccTE=?C:B
.([d<D]_2baaI54VU(9_W#O[Y<bHS[#2P3Y=A-S7);SXb>NW,&-gJE8J=3/>&7M?
PLX@YZ#FfR:dQ&TV\H9]_8&[G9OXA_bPf5QI_Sb5F+>CB:YKPQ5)0L\)g81W)QYb
e@;3<[]Cd7.a#>-1#C8BabYAZ@gH(8SRQ\+JP<BS=EfV-)4.G(<4=OGF0V/90\:0
^D?8;CXM9XPfT.?CHD9B-\DA)+]0>?318d#>g09]4D&WC84AgHEd;(&#[6eZ24]/
A:aW=7JJe?6+TXH1^&CXVW0-J2,:A4deQ_D4->OHe7<I#^N@^CJ+W]P6#fBfM[gZ
-1_5;Q+EE.29XI/H?>gGf:L;fQ6A63_>M61M=N1PeLK/(=-?GIVM\;(a-5^3<3,S
RFgEF#^CBYC:;QC)(6#QK9_c1SN.T/>;dC(]N?Q3\aY[0<(F^TOM2)&d6E7^UL8-
A7&3)aDZH1_L]^STZd:ZJ2[0QL7Cdc_HMWQ:W;PL]);(S+/[WPbJa?@)N(L^/[/B
T&L.PDC=7X6J9@ZU,D/c6eb?^\eSd6]b@-:c[\R4Xf,c;U.;N/FB;#UD<R2>3fRe
JUP7Y]?RO+#+A>\RdS1S@OB^C96?9P^/UWMZgUa=HC]3D&g16(S_KWK0Oe^;KN?S
N,/H)1FfF(d5<)2cD]VQP3PA8&EG2e)#3f.UOZb1DC7@^\bV=g?.VIc[GGc(J2T?
:)KeF0&YJ/3KR?GC)C(PZ,dKIC7.;@J&X<e5#_?d_:5M;[GLR]HDW[AL+Z2Qg>:d
;Q65?(5WC]dRV,WJRE:;EW5g?gI\dX^,[adV9faJSMe8E^;dJ/1g9RY#,?>a^^H&
I5]Y/0C4gX(,<RA1K\)&UI+PK[=G&QLJfS8K=e+\VG-?X>3dW@Tg-EDPg([9_b=<
TF)fLR23CLI=#V=;<K,c3F[PV_3+@64?=f2Z_D#1L+:@#L#Pc9Z4XRMdCNEE<&(S
I0K2=ND@)eaW1(e[]I_MUH>?DBZK.#T8F),6/L:Q2#1=^2-)/cD<+0[447[@4XL7
AgRLSQ-cN;+JQUC28[e\51K6P9E&+:+M8HbJ\aOSW(:HBf;QPS<(^Ia;U35NL4))
#00O#.2+>/^6KeM@4E>b.#)0G;E]V:8],&aCA+Z)^[(3SYC?1-[S67)7S<UI:4R2
JX::A^JA94>_Q@2KTCZV&B9cETVDRM2&\[^@BXaTH9;,a:IPK4^QYX83]M8M.C+P
/?2A=J01#^Q;Q8YK+F6QE^?04W2&3QVVCgJ:+LP76J3(ZPJYf\d3QaN_G[[I]WS;
_VHRX:A7?O4]<e0-BVESQJ5^<\cFAg9+=Pa[@5\BA1a[F;&@[9eHN+H7-B],UROF
+_A5_e^&NICZFQ6);YK01@=]3W4O#EQD115dWbVI[WeI>E^XdXH>[7&HB;\-8e:=
02\(9E=,V8JG+Y]/dW/V^YWK^#./a)PM1VGSN#Pa#eO<8_76g1P&2I+^CM_&NO<L
B@bJe:.dI,DZ471Da-L,&LgfS8^FG?2UZ^?KR1_2^gbK1/#-R7D#:YJ/0?M>^I3C
\]C[X/S]1@TLUF&bdc#dG=)?P_FPA)E_\_\;[5=R4XJ&db_I,]EGOQ51KT96(2Dd
I-eV,,1\X^G5a_Y9(Hd.56D3FY0[Z?9O]:/\5;8d5;V8c2(,EaL9]C8TVJVXX.a5
d79&85NY60>G(2dR?C?ID=82166KbM-]Q:GC3-BdO1D\TZTU7c;LVMU@2OX>NOO-
]42JHZdS\Oe8>;N#9UT&LJ<6Hd<;Z]Ab)PD:&_MU,Y-TD)e>T&5&3MC7-R/4;L7-
3+\.L/6[J\OM-1\^5G?M5SCM3S?79^7RUaUL/Q]W.AM/=I6>?=F2(GV->2JL355b
UTHG;-ELf4e<86Ja]7=aOcD4BPC?a.)gXUF)@LAFa_U=O_VB1C3-D+@ALI,>TQ+J
aX8,#dY(.(I0b-TaM2<[GUI@K+#YI5#eLZD;S8/V8XFDKVS)7GW;G+41C3(6??G^
ZB;_)D2I?ZGb(,U>?W9MKdO3>U,1eRGT2eF6L7J4LPVT<..Y)[]4>I#N\/@/UG79
dDELA1>fZ=6+CINKQ6Cg3[+E0YMEDgFcc(,D2HU:V/E];EN\V[R[^EP4T#Ab6fY?
#^+&HSY:,60R1U_N37eQbc-fJ9HTI(^6;.+^P0ZDG\@FS\]/+f__E)6=e8E.,QV?
G9AQ]7@L6bOAF<ROHIYd2Wf8.VLBKBKRVI_R4PA_<KX.EEZbCKPPSQ[JP6#4RVCH
<T+#X?\R:.O,CcRN)]&)R##O@OWd=,HU80PFKGfI>ea/NV(DM+>W-],+?<f;XKYb
#g(VG\)AN^SNbBZe0I#<>-8)X)Z/\)UB1OGJFc\BI#/C25M@=;<K_KI-O@N><]D5
#+\S:WW:/5I1([)J<?[O)&I>CR^N9SEINJbPC[gB825#<b1S(e_^R[;RVKa1@XGI
M1QQfB(7JZF@ONO0>^HGF#F.gd1IJ-N>XWPK,7ZXA;.?NX5fG;7(G8Y:53&8Z^59
-BCf\DL:.g\a[>JCaMH<CBC8F<+LK+S.854)?Lg-@2ZE]O&If>7gHM?\60Qe+\2A
Gd@=cQ#8gd4NG\gJPDIX,K9E@fM296++)J9&7Dd=,WI[>I<?K6MQAeYK0c(EER#;
9He4U>WG&KH(2WORV3Tcg^>J4aE9]8,X.-7e=Z3&13e\<1M/27cJ7LXaE_P=^63(
ZgDRI:W\DJ[DSSJ50SD-fM]-6e1Q_Y_0/(BER_2?2Ya?g<7SO,;I]2G[-GKY@dZY
c0_HH+Fe&_ZYe7^DG/Z^[OI=>5\H9N4^7VLLB0L^=;E[-C3YC]M>HF+G>UGbKfc9
acMc)eDVFEH.@#egd_#?+;D:WgI</;DK&R;SFI_7<fA(.JSV^>==Sa5XI&QJ4QIc
L\&:G\X;<=W5T+U+b:XVWe<c6/X_[+SMd)O8)/R8WK,6C\\C[Ka+b2O7#a=@^A=?
WV;CLb)590b/38cWYD](:Q1JL-Cb4C\=eT=)&T?AGV6c:=;+cW@F7fB&CAJRVE;;
VAW1faG^<TWdMASPI^?DZHQ0>aAaI]KS^4cX(U;#RfJPf=Ue#[TB+SY\_V-2]JJ5
BRVN@;\MWPZ>&V)WVTd)1<S9Y-B4)@g#:#</]E3>a6EEFPCA?B7KP5^D(:QgdWUA
8XX>T@#=IG_[X3<<+:DG03G;0\Y_,Ec-5AN:HQ]7YL_d8O\+]ASRWX1N+HS6c^?E
DHU2M@4.+#D8C/\4;P7=9R[9cV,Y>,((MBS[/Xf^5f-2OVb;[-g]#4WbE[40.Y72
]H)TWE2bCKU]B96^M0@KP:7\QOUJM^3\]GG(8@Q2W\3SQ:38SVbS>)8R\g+RH<+V
B-_)GL+]30WQC=I@gF2aHfMK:E:51g5M[REWC98K4]>CNbMNa@[9,1S?Z2YN.bNV
L:TH^1gK3VP5@@__@/.T]@a32^K)9cWRXCA?IH53]NeYZDOB5\V\]4T?.N=-Q8>X
=QS&4&;Ze)315@S>;6HZ#=R/D2(/84^O=#1]G7>0)8XY4>+0-A&#1Q;>-L1He/Yf
\9-I))9]IQ@8/P<>OCa2(1YHR.1aE,]K1#VeNZ5GY,/@)_,1dD336IQbVP:Z>YJJ
DdacK:37IT9dX#7d<W&Q78#>0=GNEMYGND(3d5>,(K2?N5[T(AD:[:M-@f(<4J;K
0e;5ZSeOA(&K6IRB.+H1X9)?bP0A;,N>8V&;?FUR=?H)DRd>.6.LG<+G&@)0T\\-
)OF>A_PEeZcYZB[7T3RU43BdbE78VAAQ\67Y;T]@g>S_CH+BDMf;EC-(T(9=ZR4_
D[W:0=N&=Ib#.UKDeJ-W+E0_4L].>3/^H<:D@F62bE?f#+JP2M3Q],0ZP]\O@gKX
=AK5Q6..)59\2I<]^IRVAcHOQX[S9Q(YGZ33_VW@],2X_Bb3FYK0JM7g^a0eM>;b
_F42Z9c&\R7-R1J/YeHA,G)/HGJHUgNLe5W3/MZ8NQaK+BB4eX[aC[6OQ9K+D3]g
#eb]BL#&@#T:V.Fe6VSa?(1?A/]gfJ2_&_.(M1<7X\46K.fcRJ^@E92#b&;<Fe>X
gHMF;_I.a4(#RXf2S[)RVVU7;fQc.]9UIL6;4C)?K&#/VR<CYRba+@RUAa:,]3[L
R?H,4#0eSS5J+6g@&IP/;8&+/@#0XEO=B\c3>^X&C386\a?4Y]I&A>NU=+32@<ZY
c^UFJZ91E@7L/.>aD;E;FPSV\&R5-[/S3g,0[UPacYO-MR+UV:(RS:d<R8U75-YU
<-/>V@Y&\X6CgXPG4^TU1PMUe(TU,ANU1^@DG,JO0df<<HJa\D_81:-ObPJ.D]d_
6G1&2IQNc2Y,>dNN+:G#EKAEgPRT=WC.J]TKP0(<P]S[)&2H^<L:[Tf1fOgSJOdW
)Wc9)gb@?(6X-Q=-TG,@BTF46]:8XTRNBe&MQV0E^\ME1/AT#45CCa=ReFNGA3bf
PM=X1Ja+e6L\c?[?QT?.Q<eUGfa>:JYL[.#T#gK<T9F_bY8FK;6_9(9/ZGKCE5WL
0/UZ:JJ;OKI[B#-]8aY?1KED;,\1/@]J<FHa0d6JOAJ4K+(C:-[Q+UfQAZ:U8OFN
gGE@W@d^)X_VA)Jb/f??>STZ2B4OE\?g,9,>MTA<ESQ@8fY))Q(25N8d;)V4ULZY
J>cWfa+)A+WK6@:gOC=3_3KI_@+8E;[YFg<1OA4e/04&IB8)I3EL3G-DH(NP6SXD
^\@K&X1Sb@HFK[U_LC.5Y1<BU=0T/;GR#S5VGJ5g9-:\:\?4,D-Tg=B6L).H(4DI
8W<e(\K?Icb-;ZX[I^;Y,00U6HZ1ae7+OO=;AdES#OE\W[aADFD9JIaJZ9;@U,db
-]e=G[E)+^4/H)e8?d#YI.??UG>5-eCOO@U15VJ[>@<[W(\K@5^fc_,9>R(OL[OP
3V;;UHU;R)F#AUcKO5;VE#L./:C&Wg_GL/b5@<Y.9JP3+X4TANaYRF/G1^L8eQ?[
P/.2HEP@NDOM)7G/B&60))Q4ef,3:<:[T:fOB6c@N1/AOVR#7M)HH@S\5L.=Da9;
DBSD9HRPO70U<II=PO=G>Jc]21Ub8)+0#F,SR&#ON,aU.CKX]I[g245YYQ]NC@CH
e>RcZbP@]]4I9dGX7.4/8W,#A3)^97PR33:CLZDX2G1V;,ZaDOEe0>OL?-0I,+.R
&c_OGPfKG=PIV].1\/+E^PS>NZM;9BYbZO@5SAG^M9JA([AZUg7TM_&/D4&<eBRB
6Ee80IAU\d+KLfM<G9L)(]b0eX=_9ION7dAA+C:0E;C_c))&C\BPfQVG;0dES<#_
<N-:?&OOTfP<H4cD<5AM[OC=Qd/8bE@)M[IK<@<E+MMHKZ&G-#<X4MV;JD\OC)7U
&BFRIb;P:TTedCNW4-,+6XE2L/]fVA<cg23_a]TNJ9c+DP>=G2&BfCQ?H5VC,XJ6
.g>YgGOME;:#U&ZYaF>3PCX0KXOEaH7QgOEWa5Q\)6/T]g8M<&@Xg+_1EV-=8HX:
GGSA]>adR;N_95;C6+Yf\.Z[W+IQ1[eeJ3Y5SOH4DZDOXEc2JMP<6Va+GcF<DR.[
g0.LA1(&6Ka_,O5,2aUW<I&NYSB@RL:a@.,/P4<eK0d;2(5a&COR/c^LV&1;4SET
A_0E6.DY-I,H.0/cbc+_Y4UI=&Xa7aLJ<,LWeN_Aeg5#A>+SBH0@<-/UJ5<94H7/
<GWJ+_CVX:UGRR_\S8fTVWL_RCGV=[R3@&OM#VNaKD@eZ^0VXNKQXcG9L64-9\aU
7U9XYH6Z?=Z+I[ME(;8)SQX<\ZZdFZQQ7D)B;Z=f0aA>FVQ^b6QYL]CXI2b7(QTd
>6eV6]K@9?<HM;&Q#OAddaF+d8fR88_H(\YEd^,3)5GC?:gC9ONJZKWS/2ZO5Gab
V-/GF1L^JPCFNDF)B\.eX-f6SR08f.IM1W00RDg3LHRZ4MaaF?:DHT(B\,SM&A+0
-UF#f1,4SU4_(3H>(C],/O,G_SRbQ)_1+=K.CZX4[b/V5\EU\?.XTMJAa#O6e03@
dC+8KgT(HeT1>@0K>9c8QKB#L)4Y/-LKPNde#&S260Z7e1L.H+&beO:a\g<J@8C>
<<?BHE0+6/+DU5@3g8M78[fBJ]1GJ;_UE-eB1A7Y,T>H5>.@MU:J9=,[]X#AR,6P
70VfCHWFd9M^-IM\>@,,gNECN0&dC@^bg^e2@S@C>b)XPJNRI<PIUCG=DW7K^gR]
@=S#&VE?V\d0?:J#]CTRaIDV5D4&JI87Rd=^Z&\7d/4Z:TQR<Q7H)8.-HQ.8e>OA
?F,-5N<);P^)JTZ?PeD>69-NeKW5[Y5VJP3+NX(4IXZUD#4X&cFSW9]Y1:R\VO=F
b]_<e,:<RG74N.dCQa?cTJDT.&Tg+;#-&aYTHDHI>7PFCbf=YZ:2IFbG83eR#Y.Q
KHO\S5.UE]K+2@B?db:(aQXg?L8DD57UJg&&FLH;eAZ6#DHXf.6MbZIQJ6^5JN6[
15a&G(=dO:(MV,A,F#OP4T;S-bNUMR1Fa7S5dX]QXJ_>[3M29@,W5@(AO@\YdI;R
bg^>C0X<159V)g;.(464-/3(;+60c[KD\K-M]-LH6PYTfF(4bK_;-;M&Ac52F-)F
1<1f+DVD>S\1/LC.CGZPW+QCG_QZdg(R:Z<TUW5ZC)M<7-O/aW\M-3Y\V5cPTd8I
V9C/bP++1]=IZK>[,F^;#CSF3IRd=bRG#e2AH(?S&I(GeLJ2MZDH0SXX34aHQQ)>
1M\9g?:JH0(_RTGX(V80H]I<G1JBJg:e8VY9PeUX06fNX@)3/XgL(I3O1;KAM&>g
Be&]Hg,4A(fR3N7:[bR80#c>-@QDR-]+,eWQb?L/)QdQY1\A;49Y6O9cC5/L)],9
55Y&(:+[f/S]B#48>.M128@dE\-+X+0E.#AU1^3\),aYBU3XTfR3;A5Wb4ZW@,RU
QZL##GQ0C6;Lc=T./EYZ#S<14)Da)/)+0<9NMf+3]&UDK&G:)M@&7^F09P:5Gb\+
D4aKDdIVDKR.E6SZdgU?#;IS_#Z;V_BCCPeIUE>Q]^Xd=CI>9cd,ES+OB_HYQgcR
(Y3dQX_.J3fDO]@C\8(5(=/6\^eY78XeS7._T&=8?81;V]8V)#1_AUOd82SbEe>\
.bebZ(@[?9^GU5<+7Xf994>I9FS?[GF]e#K#ZQdOe9?PYEHBeX2OG?QKAeEGX90[
8:V4XecR8?0ac.2-8^Y:PSfa0)H=aG&@@9bJ?O,-fcGZ(S6?,F+XIf=&]Y0_>A3K
^4fK?N-8-e=^1=L#[JA4_V[N_>LO;.[Z./=9_NeY<fWY4.CP;<FK#4H-F4eZeL/&
U9FPfLS)OG#UM26/C]LYN2gA1\-Pe,B[EV]G#=,b<X_9=R1aUZUcA4_U9HRH=<\A
L&4H2da_e.:_NUG;YWE;Gf#1U(f9J#/J,,-Qf,^=M=I5[MA??NAJdLMGF81WU>PV
_ZS?(Z=KIcWVTf0FY26(4cO=9GFYL3Z^ES>H95S<BZI8,g#Nd3)+98:SE6>:9B^3
_)HBe2RTf+Nb1^XRZgdb^Q+VZ@_8c#]U2Q.)[OZ0[-_T?d\g6\M?8F8+XE4Y63[0
PRU1GT+H,C1HV]Tb4D_.C-_2Z\W276-SN<ZBd&8]7&34UJY#W7=WY5=W#EO2K@g]
CCD=cdN2,V1]N2?.TB9CTSdK;e\<)NO//LSSb5F\5d8<3?=[N:eHQ.U\L/&,U\c?
ab,Y+A@gEL2=5ALC9?=:A8#8),+R+]N>^@)^7^N@\U&ZI725EH(XT:D&]7]U\FeE
?L_4Q7Y^LOT.G9IG1V]3JX+.YKebB<B/E&6]3T]1Z6Y@T;.@cZ1a,0FfGXA[d_W6
]dI[UgJ-1/gEBa\<T6?KO5#Ua00)T3X\c]aTQV-OTR@J<R-.RY21M@J3]_PWHDdZ
@,c5GW<PTYXAe;=K^+V=@#ZHSTX-11F,54I2+99\1bSW:&9SSCCZDD6=O_#\NNIW
[C4gV08d:UR3c_Y/+[>&cc-A]CYKcV1MP)U^NVK^D14O&fdCR.,b0K-e6R\Zd)6\
[#W^\5A1Q?SFM/dNU\>]-0YBbMZ/__ET:b/;ZKa&(D+UB7=[;3KbR2#G<dJSTR5U
(Ob#4^,Z5:E.F=A7W-d+]7/87H_;Y,RfFaFfgg^7SKV4@TT.B+b+2W[)(:2=cGO+
2Y)[(Ca-_G&?NQZa/1cC.QNg[E>RF>V/1?3DLeWL1WADJf\V4e,dGSEc),aG_\O>
ID:MQ/ES&JR/MQ1(IULG>6:4<6S&^-FD]M\\?@;gWI2(R=b.@U\_=6)@SADa=3\<
DE@L,dSA(F-\6<9B<H3,.5&bR/6_3b0cH]),bX),/,TVI&3+]>W1U4dU)KW815U-
c>@-DNeC/0?3If\60=bQY)P#U5OLOLJ\c,-cFSFgc97,I55>?)gQSICH/0fB6W,@
Vb.aIO>@/,)2Z0D@[/_DcS_OH>+aU1.0ZM=4,5H3]\6D8IJ_)6cN5B^+K:\</J@g
7-]>?WXXYF-VO/(L?D?(6gG(K/a)5\Z-<.[eMMSMR,]:A3<e<KLHNCaA:Pb_Z97X
&0Z&N(5fO#D9Se0G6/R^>-D2@IYMa[5d0O5bb3Ng@[@V\b3)cCW5@CZR_6^\L1Pf
FW6DGT8R?0&&<S@5eB&K&2;MP)(M@_=0.66db)W?>(00g.4H0b7R(1K\2XF+KJE6
-:ZdPB27HeW+U(L@0F8Pe=C<#>Y=C9G/dZ_VS57O=(7M65I^GcKWE/X6=cU;BBUc
)-)Yg.T<T(G_SWaRY0F/57(:9DOM1DQ.J98&FK3ULMcPaEO@:cYDWLT,d[[1b[4\
0/6>>dPJdaV2X#2S_c1W>7b;ZcDD(I9,&QMYQ6LT]YF(_Y]e3Y5K-?@+&.;DI8PH
SO-W8,4/(L_OYa8WV4D1.N&21-\WVIPb.8^a-g\N:XWF</f&KY)B>1Zf/>eQ4&+:
6[UJd#U_dKBHU-=TM=f<bK#<C4SGA?/+DZBIYX@:(e&?LK/7^b_(P[3\Y075WUAT
cCc2M:X,]D2-Y[5\4UZ>ZcQS@38V/1U@U+a9I]MN.Ia1VE+LCI;/&06Uc<8(?ZHV
DT&H]+GD57&^\,DG:&8.V5[1H)@YK+1:a,\T;T@g+3#;X/O7D+;e3UX-/Lg5BCg:
\AcMCLRX<HMR<cDH6.JH,CEY[?_/9ZU7Le2I,d8<2Qf0b2W^[PbF56270IHGZMDG
:.)2AJZ<UT)-FU&JL&[Ff?_Q@]L]>BX_?#6[&RH5+TMf==[O<ZT:JK&BC5[g+8cd
-\a8DV-+X<6<.8Ae,\ZRZ=Z=.CHJLHG;fOeYAV5f_b)N3<8B#aLJU;#-A5KQeY-2
D<cAF6Ce&=MJ_,gE.<P3^M:/<[Y6XAG2EZSHXf,VW<0_\T6P3J&^O:N:^<d(Z;3d
T5/@e54=9:]:E0I>aM&.?Y5_0H()gNNV=_#)J5/FZO#S;aXR@YXUW+KN@?L9b_Vf
LfU?M]M_ccWG?5RZgFMe=)Af&0A.#;X]]<+dC=^L+E+(UJ^&/UG_ER&0cPJWfKeL
58;Q8J9VW7b[O6RDKfG62_PWbg/TGY>0Lf29c#3GH-VE0B0:GO@=ZAK_WX3PZbCR
][LLB:<Q9EcQd<#H6&1gTA5dF6dY?55HS4]HF6e_5#&.@&;Bc]W^AA7fXGLcd[5,
5:Q7L_WY&H7c14CRWUN9b4K.2=PCN;8:IX[M,(2]ZNQYCFM.A^F4WK1+-Z((Y57b
5DB7/-,/aPCSMQF6+@9Q,4dOaS3YReF>Ab,Ob.PKAS34Ye[112fbJ,dgSN]VW^QW
=]/;c99]EK>S1OLTLTQEfP-;_25Ab#8S7(._50FL,<Z1<XPd]]]2(bB9/JSMM2b5
Da5#)^@J]=?F3AZ9:MAQ_YDK:6>K0-7d&<.gA]4-_bSM35g65I0KYUQ.GKP:AZUT
5<8,0&(AFCf8:AB@3b(19d]?U35G#;DLGc]D6(]]gDB&FW8;fZ5Q4QP<5=#O,\>K
8<_LEG@[bNC8RcLXdD^U&4[8&@:6Mf:W,CXFA.:J5a=F.#GIf:PIg=KW?H>>T713
FX@F#e&H)^72?1G;QIYc-1L0L-O,13@68>JW.N[^VdG=5H8.e1=8Ka>H8POEC@K_
a)&)Y\\9TfZJ=?^YG+cV+g\MeO&X.PYdNYHBcNO8&F2VT>2V.a#ea04NKI.LgP0N
fA/E&+/HTN5WMW.?b(W66B2);;VX6H=b=)004MH.]FGa0(4&-dO0bZae72__dG#I
XZPD:)44XT9edR6,3g5Y>6,9aE-1bB3/9TT;O>W\_D,0DBX\cDM6JT;QKW<TYP>S
b4^G\774\&@^+++=dMF7)[@c[)d[/WN3W3bUc?L^9=<=Pa3AKJbBa62a#B3L&>K9
YFBU;D+H5;@7fNWA0+DgLJ?YKRVP9ZUaV)K#O:5<[79/BNA?:aR=Kf3YCYU]]9P)
=d^]RUB9:YTDNB:7N0-eLIPZ6[5,.aEcd4X0BgL-WZU=LYZ#U3Q_NS^RY-2,SZ#:
WSZ<4P7/^R(9:E[5VQ-P1a?@,7<,>aAV9U\I.&\,N4=0Y>FWN/gd^N-IaNSBM9Y=
d:;?:GAPP>F0cRA>ZV]ObZcI.ECVR^_+0=H_E[+O/<ZK.fZB_CDQ4C9Q8RfJE]GO
4beA=5bMdY^]#EW]NBBR/#RZ>;@)\cT3P\fV5gI;ZKDbJMQ/RWe3cH(/)2IA]/N^
^IDP?a[E;ZaHcJ4=:0<<+Gf&@I<FZFSe:6)P7:>GY;M5Z_2;754)[#S6S+d(?&U)
Xd\b0eI6cX.X<N<JP@7GM,]FaV<:S^dBNXHTIN.,5DfA#]cIaHDBPbAUJ/N,dV=>
[&3/OJ<a_8e/[:d0,aF5XZM)?GMK)])gRL&48KZ=Q?5-T__c,Tb[;_]4X>RX(&cF
\>ZWHc,1WFNAc1b9QN-0EO[<Z@6J[b9NR3YFaOX4NCDXb-.IE,OQBa,2,^\7]A;b
D50PMF2/eCAYD#43RgEESSM[JBbV6bCb;=<6=UJHaF+#@;9g7G?H<N&JXR5^b&&[
EZ&6&D5JcS]R-Y/YUc+;]D4UA<GLY/0K]3X\^L?(0_C]Ld3MP#8-5:7AYQP^YY1c
ALPS&0BWaF+bVGG.UdYFYYV35Q#.ZWBA4LfI&<V7#AT<ZB<g/8^BM+@4D.B00QI;
2CKJSb+ZN+5[H_+_3X6.\O;+a<ZU.Y8f\LQMdMWQ3=Ugg6/dQNY0WF@<Adf0-eRL
?.dCSDTOgYF+g]:ZUGGZU&c8/K<eLfLQJX[DH[9&LAXEX6O&c)_,,1fBf/=+K-&Q
<O<D8R9Ee3HWLXI[;0H@g#&QBGf9e8O@N+?6D4/J^/V_9_#G[K9=N,]IdN6\_RF9
.IaO0I8;)NLE&Z^.S5S2Y:LU3,E\e0A&P)MJba1gK@).Bdc-S5Da1a<09).GT3>9
_M3C[Y:0.TV>3)b=5=Y-e/aB\8[IbB=D=4H=f5-AUW44]8O]_9=DDWDK:0BFY:AH
(4ZM:8]026)SBS(3DD4&d#.EU]+Lg?@b5#a9b7e]6@LW]5-I;0W:QG=AB&&B1D#,
Mg[4<]=QGY(0EUE><1X6HMEE4[FGNYE#ec/+^?KE-]Y12:TH^M&dN3;OFM#bcc\7
T^T,VW@3,O\B,^]7#ZZBPb##IU0(cBV0X8/>,.U4DGVReRK-VWACFN23KUD#-:J<
cLM?TA9d+<=[d]<,?-+KAL.6Ab;Y]L[O-7DCb.CNWX-=AXTf]Oec2PZPHOO3A&:a
]>P>QN\/]LJ\&CRLOCJ6EYH@bXZ;84;RB9PO@^0dQ\;B9BOW[S-BCCd5RH9/c0+U
V9Y4@F.=5ZcT5@0#Xc/M6UX<4_.g_MAJKFW?G9_E2U)64USNeP@/VN8.0EXCSX>^
_]E=T,B3XO)HabK1Rg[d@HGQCc7B#=3(^1MU8C3V)^f>6f11/_9@BF4JQY9d2XU+
3<f]^Hg]_]SBPUc+WYdFW3\d\:U9&W4MOI.P;KbZ3YR[,[\D[g?:K>V3O#^U\Tb&
V6Y?/A#(g)R<8L(7O76GFNL:1Ab@1^W1J?(,De]HZ+_&(I2<6:(IV3E3SOKP)AdU
VS(R6,B5V=OaASW+N20^cG(_=L.dgUaJYRY[7N65R?PX3&b,Xa+e[T.WA?X28g&_
Z<7/[QA7H7gcB:ZIb?K>&ZYAH-..Q;=^#QQ4bg/.M/<7dF9&ge<(BRTTT+Y(fC,X
>+]d6d^?\H5ZS(N9:B>)>\RRCO<<][F&)aXH#8[]]@IM?CWD,WJTV33\(5J-&&-a
_7];RJ&ceT0I9C?7I?/@;#L)#+7X++M<S_XA)eO[HQQFS-cX?NU=YN5Z6EO?.#QN
A5_Jc8>>b]L7g.C4Uf+HXA7/S<Yf]XK(05O/WeLPED4/\.&BcKe,75J>fCLf._^7
3)g<D-Y3+]=CCV]A(L_T]1HAP9V9^WE[2-b1PGd1;<F3<e1RaZ<3/cc-(07g<63M
)8@=>5N96O4RY2R>-0T;cFg^&JgMF:IT&2VFFG&Ab]U@M=SJIb9LN]&CK]=7^A]>
gL4/>-YIVO[W:4(X1&bE4W(?SLU8+d./1DGHYBUHKEMLDaN]fXc4OF3M]fdbHBD3
75JQ)HJ=Y7(7aaYPWX4[Mb;(:NA:RFE2#(XI[fR:947BG6B6>)\ZL1Cg[:;4EHE2
9FWeJ#C0[;9C?+ZC6OVY7ND.e)Me_@#X?E7+_:CB6RHc<@2eMM)g1CJ:-d2\J_C&
TOC1D_.Ue-f:FMV4I2bg9S_RR-Ka=9778&:MIcI0FEXLJaBVFe6DZH37aDI^1H(_
56#D6JMgC,_@1W6X[ECD5:?1[BEL+FcNP6UX3A4H,2XIH:/61^S)M#<F49Zg/fB)
=5Cb?+D9U/Jd+A^[D[FD(X.K8D1-3_TQEf^816II@H?HbHGKb+)(6:FG#NcW/<,D
^>E@+ZVMPC3A#)J8)J(IM,O3F:1F6DR-_2<<?DZWU&&;8)fVf]C.\Q[]2FLS<.[)
Y_:ReW9c4fF<7cTGFMLRA=7cC8E+;S9FVV++LT8B57DKP?60T[IdV]VX(+YSO;BR
[3K]V.EL\9;FU@H55L?c5>C2.]VE8:1<.Pb1?YdJ=NF\TGP+eKO8bfKgfN/Ub4=0
U3Yb1C.XN8EI?Z^<BJJbK-ES=&DKabfaL^O]#0bfd[]GAO;+dU[^;dWD8&QOX]Yf
HT?FbXDf4V0O)[bTeUEEG;&,+#T84cU<17=<L#a[Q2a>\;1=VEgC)HL+L-,Qcfd9
b(bR8,V@E&8HK2H0H2_Xdc4U[UIS4c.;+UM=]3TONF5eZOW.&Ug;RBeI>:3K[a7=
_P?5IaM2KOP]BC^[-F\3(D,A2JMO\@0bdT]R#HV:7N[JJ>,4]R.I=L-<522>4X#D
^f3(S\g)N]KLUJ.6RHg-@N[AAY]G)8B&TgU@Pe50)c;=.JLWXX;JUU>:fB]U.FgV
?8_[2W\V6b\=B+NVM]#:b3#006>?JN8S&YAA#e<[EFYe^?H6+]0EWL05/WEbTJe?
Fe\UA9RVY4G.5],;4f6..:V_Rc+2,8Z0JKMN@aO&3@8GBdD?cEUSZ/)I20C1Y?EW
W4C):Wc)4MD^72Ee53;F99eA.>d4]6B=9MGDeLA>b5gXA?]T40)b;OeDYF0^_?SF
g;/T[[O]H)8Y_3ZW31(@.I8ZT<BB8A<S2/9bF1-]5A&bZ(A@3S^Wa\BdEKDgf[=7
ORa/S:CX2@d[;gQO+f(=gBU0/[,2.JD@;a?If2a9W]>#915RQ,OY0_:G[@OTU&Ua
fH-Z;LMN<DHMK1WU__a4-Ig??Q3^AD,J8&&a/>N2e/03.HHQ\1<]B4^=[#6R4JG#
M@-?&M;RE9:cZ#Ob78X2H:9c<a&)I1aLFFAVY9,CeM<PXFF(@ID+1?8F(I2aZG)<
GJTE/1PJ<g>89LAG3SaeS<7=PYc4WWf-K]24NZc,aHLM>e1VD0\@DC#c.EVgJRLH
YK6fWKAf)LEGbG@K^?Z?4FM4#Z=X1b,[2TUC/2PRC/0;42fIH02EBW12Z#eL465G
N:4@RP<X1](:\SaG2RVN_M:\7I1?^KV^CPg.^V_MJ9[^#fJG=FJZ[0/0680&OJPZ
)5KL_=3^4E[@Eg+18Nf>[C][:4I#B(65:\AH.I;HafM7.T&VOTV.32F.+dD.O,g<
JB?P+W/B?MH5cfC3LJM&7Y_??eg1f,5Wc./E(_T8cOQJ?7GT1AQ)FK\H.G+LaL3&
8XMZO\[#+S#Z+9J<HU<G&&^I(L160;XbLQWA.PReN8b]ePfP1@>-I0Sc+359Q5M.
+C05J2Uc&QN/4JAb=.EI7_Fbce(1gH?RQ5XGM8c(@QXcIYYT(6&A^R5\T;Xc7P8&
g]SRCWIZ0>88@bbWc3Q2U>NM(U3=SN(]6<Q,NJC^^Y+bC6_9N?GVK/VN,b8_e?9S
,</DU[/5dbeH08TU#QC#W3BUFSg\5^cN<KH_3d&T9fN(JSUCHY+XP]D#[;<;HHWN
\UMQJ/:Z//0WF;Y:QV9360b:WV5D>SbdgE[XEO,.?H7@G).G,6=GEXNXMF(W1/;3
Q5;c=cAg/Hca#8/G3[;I8Q=b8];LH?O7?XRV?6\L<a)P2QMI1<SWdQS2_35[[YdE
\G)6L^5a=XYAbfO8B,TX3]&#249dTcJgcb;.>gDUTBd@BJ0?#NO;GOYbI5J#>IPe
KF+3_S7/1GY;c-;RSXUfS+N8(C0+>=aC>39[&KI/9a24ga?MCc;+2P#g.8BG77<[
,?\KK&AF3/bX_X<dM168AO>^gF;A>T:SbJ/N)DI&ab,91&@1Z.T.f)9dWP&?NR>g
I\GVA8C8([Ld-Ge_^(E3S@a@:Efc.P>aSc0WZcVY>e]G+dW+gg^^JZ-PEcf3\\4K
ae5e.C<U7?#LMJQ3e,2b[&[WK<=BF4adEg?4YZP^bD_-=Z+XK4_5SH[.E)fgQ[Ye
f:Lc(Y52-OX>84:=Y)X\0af4gP@[A?-P8f+Ja/bGdaRQ/W(BTU&&\[9VT4.1-@H9
g32IAQaB<85d@_-EXJf6_g,UBRYK^4d)VI4LG]c0C^Ta&PAOK;]P=FeJ(aUM(c20
2<VE1=/4K/+_.=<.,\#BW#^C9&#I4KVLU1\0RCIb_Pd6^@d+9Q6^95/;b)3/RO;f
c&bNAA<WN#MHHN4XM#Y#PNeI3U8F&Gb6K#6?O6M]3C^@48.BZ^R7@A3@R&.D/\MV
F8TR>]Y7Y.=9M;:AL@1N:K]a5U6Ud/Y;D6_5#YW;3ScYR&WNP2\@a5/;XRdMTOI+
S<\4^HFM,+U1GAeV0(G9<XfSbM^IDIPX-QY[7H:G4P=O7Sg><OJ3U5#WQ)g-Df1U
g7L/0I^E+C3dTV^69Y(?c;GAV>&9Z,\025A.H]?C>4VW:/C>e4VE/_-fGZNL4C&e
6-RKaTQF9L8TR1bTEe3Xd#5[2OTVc/bK,W.GaYOggJ)HgIB2CN2YI\QG/b,_(@@-
F0AA+5bU+R52<fU0QG)^/5.V;M<R-,IcM1^N#,<RfWF/])aPW.GaJPJeR)&GZ6;(
>9K7]\aIBJBUUdfFbB^Qd-7_XH1+&+7.Q:XPBg3ZRJT7fR1+V-Jf45@GaT6aeaTJ
\6:3;>)4gX287SQcYOKAY<C_KS0+Y<CO@[=K#J9]J&_TS(U1AD9;O)gI7QXR8FG.
[&_2Y:VK/H1dQ-&22DfLU_8PV)e1?fCf[)c#FQc76+^ZIdAH?J?I?e<IS8[BC_KA
@8-TNE+;g;B(?[,_P3/EL_ZH/<UdX5;U(?YTf)^(N[?eSTNF\]#)Z,G_Q]OVf1MR
XVf#./e8<)81WD=2L+82>(H-ef>@KURbP&T_:bZ1<.T\EM;X7P-/A1IENaOB<_G]
5R/W6J,[\IDA<F^4XN-DXYS,0f^^_I0?0;3XP#H=OBdS]GKSgSRfFAPM>>gM>2e-
<GHKBO-S+Ua;<MV+Z=+IC5d?RV9R#=I:6Z<L&68GGKAg<#TUYXF6]7IS_LJbSD=7
#Y5IV#@X)([2B=Q/[ZYcTVfD?;J;G<:(HFM(N#PBa1>,H[32g#\R(=A^@C#3fW?9
dCfRHSK2C6_FW@SS9K@eM&b=AN3M_8SA);&J1]3OG,cR?/029OcCd]gg^:AS=&1N
6#/e#<FB+[S3YL0.(>\?=G:O)C7[]/NCDf9TdTfL.OET_,WMcA2EBb.L1_aAR]@^
;?JVf;^6J^Lb6EF)N9_8PY#dE]Sd,@Y<HQN33L2R_,5&DW)TfE-:]7P,,ANA@SL-
3]1)HfG\Qg\#63?(2gL?Eb_F2^\GUaRbfS9&@e[BDb1A1Ig+NE4CGT2Jf=L<>-JT
&(Z:RS5/V/FJ0bIQY3V/,(9B[AM5BM<:Kg[:;WN[AR:QfcU+QP[KZD1N^[3b<@.L
[0aSZ8Mf(9GO0cWS2d&F.X&YX#EdA0&C?fcD41)[70,2\@1T#U:MVaX7-SPVNc<E
X3?gPS6X?:fZ+bDJ36f6)YPB9[\SLMTD(bL]ZFM1H(e]G<<b4O&TH?&XWOEJ-[Mf
(GKAIQW<3>5O0Z=>FQM.]g+0Ka8G+Z=_/PGP7L@<,A50]KO-8;)X^S_=8P&^b_3-
UZQ67^Y)@Ga1d89]fE76WP320>I.(>2+MbK5bA/Pe[L@7B6X;^bf7U,85]9(?aVf
OHX6G.=VMf33/?Sf7\g=B22@M5/8>8O/K4)58H,DLag5R8=G5f[g>]N^/M)DR](.
XR#3\b:RJ)b3K>DBe8#aF8T<,g(BbP3]@]>?[RF748&(+\7P5T9\Fg]-VHYK[cN)
]Rfd9]HD49:g6@;N4G<;1:T^cOcXY8B0L6e2H_+-4^2QLW&eK[f=Z;WA)^4O_,,Z
e).C0G<@\Sc?OeLG^<3(gT)/F0GDb\1Ib4_R.EO9WUQQ-_Bf5b_KT0?UR8+\ISKX
A,XFF5B3KSKUE#/:1f/B]FDR#?O1_@S4&L]W##gg<8LZcM,6G+9_\..];3H#53RS
0;VP_aGTG8&4_WQ68CNI:BY\,P(B&b<A78gQ89,TQI60JJ\(eS/PO0+c^/9<M9Se
F=\#,B29#fJPG]5Ng9WS.dS<BdPAZ4e3bOYZ=Y7TE.<K_/7cQ+Y]7#Zc^2VH:eK+
BN^UR]@Q@@fPKCJ]MUVA#C#e0T6FB&[g<gg4ZW-RUUGfAV8ILVd_D4]0FD>f/\5E
=6Uf>8B#L^7HfFbJW.<+](AD-:G5FI[#\RNf8TXU0U4X87\9R((<E:W5P[?;EMI)
?LP<ET>9a,1?4D>5BN>-E<@SP]53Y0?P.Z]a\Q;JJ:e/<c-Y7M:OE++FYS3Lf7[#
?@OT1PLX78T,UcMWQX?]>I5bSfTBFDZJ.HMMVe;AX=>+fP+0IHQbGXCK/Q_Q<&Fc
cKFCabE@X(=Aa0V;7ZP#2J0,F3;8;f7A<D@B2TSJe8b+egO4ef+9I[[f<bP;.:9K
=9.KJT:?eM64)=[6??EOMaVAD]^.PX_Bga-S,FPJ-_d5PIFG3\(710(/.8AL9@#N
c2R->HE1Q3eFXS>(D1R4=YG6/K90aS9JK)Yb6PcW,Y)H)41g.38V<.2GFX,>CU;/
<#;CLY,]_M+V7/;bN\2##>:)99SS)b/3\&P3=EL05CS([U2-H2A5?;X#0(3J^JDH
#03gJ+/HdA0]f4CG<19.6#<B9C^c#Cd1,1PS2^SH<H#TCPMG30M_4-YLS9dY&S&Y
T,0IK\Ta6a1gBSAPR:H\O+[O-RHD5]Z&;V&T)6OMSd<\&L^E\7K1#aFad^^_A^87
5a1)UMB-RNK:M9dBBVXWV#(_[FE(4=I,CJ)4?9+F[WJO7IfKPMfZAH1ePD>.8AX&
\6+a85\3#>=-gBK,YQ-#^O@[f_0HF;0e-S,^U/J0e(_#<FD=CW/,W);+X[+<fNWM
.^_J^f0;#?QJJCB+b>7gWB_Ia?5_4c(W4MT6\)>6SSZ?I^3Ceg<J0/;H^GFNe(H(
]aXTT:-@F2CFG@M]L,IJK:+^/6Yd[0.G+\SFRc7Z_E+D54_7R#N)SQHWN1_G0c\1
M+5);B5\XT;Rc-QMJ+7(dL+[9f+75B1>Z]6HO.]#E:RXgfBKOH\(/IQJUSY6MXfJ
fEQ5c9dX/4e/F]&SMJWHWEd=V\QGHA3UJd/.+TA18BeB@_TPR?:_Zb1@P,9([T1O
/D&[2/;11M@BI(40COA]A(R/BH>PL[A^\Re>8(#ON\\JSH/_R);3BbI1,U^,QU:7
3X5;J;./\eNE0R7C.Q+;=9=bRL)Wf)0F/S:^&2Q:c_#5F]4\4]I(bC76;ee\TH-@
QS/e1<d=VQH@:B;C<]YX:1EAf^9=DFE<8=]fOgO=Vd-=YId6ZMJN&CC^J^9;P=ec
c(T;4]:#4SMGV:.Fdea+cD3d3G&P/.L-[L<d/cFNMM<1O9I<E2bW_W[RDR?dIJRe
e;[:cE)ACbONPY,KI)(G5#4Z[FD0N_./>,+MXfN_M3#]7CG^KF8M;634-W@I3\1b
A][)SRNTUgWK(2);0\e([&B>/+,S]K9>6(EGI_X[a,)Ag^<O/74QeSQc1:RRJ^Y+
KgYbT]D6A]2Tg;/[RZR<D6RGQ\TBV==g2<@3N>V7<WIHQ8-<?UYd9f2S[.B52QCQ
IPAg#8^K[,P=3C585)gF8,bV0eF#59W=QR.9W&5E1>[;:P>1ZdT8,-FB(2[&EeX1
@K-?@g>-5bfIY1Z4c:2N82aK0TV[/WFN-<Ag;bQ2=+baL:#0KeM6S+<.=e^M79CW
Zg)O]G,5HE0@e^?FL?P/?J1e0a:7VRCBU+Regc>W2J[SE7aS/ORUF@5,_-DXcBUd
T+SAg#ee7HO@Q-Z:PP2aX=EZ&_N3KKB71ZE8<FI2Ya(Y0G;?WB2aZCVdaK7TE-(E
>=Y7A3[]G8[RW@g1JW8H-CRS3J<)(:Dag/S]V\?a00JbT_Jdg45e0O5:a0P)cD]2
LOZ@43<#&=dR9d8TJK9N+0b_-g2a+SPbI4VIfbGA/eZL(da@S-9TTH&cKM[_SZ7W
4F,S13T^[W=S/U3STY6a(9FdR:7LO>EJ>ORQ[P00e_UNU#6WD4[6&KZT[=@T(1e>
>cAg9A>G\bDKM]Wc?cKgG<A@8T)f[eKc,,OAZR<11/<OF2gWUJR4RFa&b8ZIYF:L
:eE/5<6#H&20R7bGaE5G@eVX6#<+>HOD@^KZVC_JZ.OGEd46T@CPMcKM,MPaGe66
QB1gP6DV&Dc:-X^ABWA>#_Dg5OCSWce0fb_:YS6=F2+)cFOU[/O>Y(5Z4J0:8D(@
YH@g967U1)d5#MDYPeCgQNcNVc/[0TNdH&^9K[LON0.UH<S2GA2(eC,)[IQbcB[&
?=)1N;>:>)+MUA&FfEcU_NFJ&V))cH[D;-R5#POa7-g_O.([D,8XS8OHeXS^g@C/
9TTP_R,Fc<GXQDaCZb^C53\>\B7V6FGQD0@M>8&L,LFJNK4V6W-Y3U0EX=?K+<L&
:8BU4=(<GDZcb@\8#++)/LLG(9VDD\IWaT=5?F)0QJ=]d?#RM[EY/)CZD;F;:Cg<
6WO\J9.J./HX>M\e]V;YW-C_c;6Y6Z4+@VE7#WU1++4AFZ<89a;JZ\L;/+IB#I_\
=3FJ[fDAfEb6eM-L27\?HR-SKYM@P6T:+S8b@L;d[EQBF\W>:dU&0U@(^]f>;OPe
A0DJ0+E#D2fSZ9R>DZ//+PXN8FRL?X4A;9&(?=/g2IZ&)CEc=<PJ_17YPT9,_1U4
8(U?Q2[W&[UJ3_V#Z8U=<cZA9S>^LBOfG>[_2FaQ&L6WMKBEb[b364J&?C<WbZ?=
Xc\K4N_McOSE(bJ[g,SOWPfVPMD5#[LUA0[X)7dQ-P0W^C1ED@d\DS46QH58H,&C
ed@;VCe3Na@,.#1P6A;XYFDH(<Ud>I(0(CDOQ]3dQM\UAG@\/LCA4F+?L2fac)?]
^Oc<A??]\).\>5M80I_bQWZPW:5EC\L=P;A1)6=YJ_KGb@<^\WgCWf9#Y#PQe86<
>3X1I61F()L.5<IH^AIC1\J0A@H>[7JW[Age2@A06e/e)79AdRHIb8ERDObR3d3d
L5+1)Z.)>H_aG94aQ6_A,.eb+g+9d.BQX?NUIIJdcOI#5CA9F=Ue>bF[J>[2OgH<
;W0JP]=g5=O/,.7^CS/3[R)2_X_ER;dQa3@36)_/W@U;&G)B6dfTB[W<+BG]BBZM
=>4=g@3C.SQ?HN,),a@[Bf5f#I=]C#13c+ZcV\K0[&HS97b<NU&.F>eH)K(0K@>b
X#V)e--eN9eFXb<QLOeZ](1W]IfE:3)Da7]WTMfFZcZ7+NaH\IM?5/^L1)d;=YCK
_I]Y=^2[G[R3-^5#:QM=Q&Z^aB/\fZY)<6T_RJ_7^0M:e,-[9\HBINVgSKVP<3TL
B.J:4NDK26V>3)PJV+5((OO./>+b=#Y+bA2JU#I;,TE)/7B9EIKSJ?3HM^FG7\FX
FEgVTeS_V@G=_=R-^.NARBJVaT].bdMCKbcPU-Q5gX_AZ-DJPGIWd1[^A^@P\&SW
AW@M@;XWU&_[FN@e=WY6Q,)<E=CA/23DT+UT-Q>:O?EIE:#YS=HAZCAB(._:96?H
4.<)B]<?8YQGFLf[:<(WS]&CIK@UNDHF-+72#=A7PW+C4&+gBe5LO<]Kb4Ka1?GL
Mb:?bN#-R]]+(M@eGKXKGbNK3M]H/U@bZ+<9]DXJ0JE6W&4gCGF])C8M1,?J>MK=
#MI;C+g/OJHN\V5)J.+dNNA?7&X+3BTd/:2^1M.1-\K#N8TF.CGEVEe1U-#DdWM\
EZP?&?W8NSLQVZWc))7,9AA)3/EHI7Zg0R8__7.7=UM)1[4JFD^)X9g^X[LfgZb?
=RdHR4YOOec[Pb&D[0SNgT)]UNab.\6VWg0(4(M/&.gK46_SSE6_#HUP@^b3c7I9
\?QG>4>/[2<Fb\UD2-E:LBX&[8O:b](MM+)K/C5;BX2)YddX+<g[fIFcb[Q@9/@R
SFT,E,d.M_U_U+A\=cZ^)0_f:0_[JV9()Nd>MDF9FMFC4Z/7F1[7b\3dc:FL>]MV
a6a9FDV@6@cP4BdLH?&RgaQJ;Jf7.UQ\A6)E_):6\._dWZ_NBbWU)_NN-?HMO/SO
]8:&,:?QH=:BBRBDYC-E(,=3.9Q<->?E^SG3]X&D7UY_C?5/CA@4<[-c8.>H_.g^
8:F&c;GcAe/1G:Kc6-+W2,J3a76L>/^CC:LPFP+8F0:Z128E8GZ>.V0YBWD5=a#d
=8FFDXF0I)O)\QEARYUA=56T(EDdeHYT^M[=1[5Y=3V,1Z+:#(6^CW/?<<0&JfC7
d[P+HE8]5WQfC1S&^Oa1/YK:LY^X&H(71gPSY.<X#fP6XRF)/7;?#<BBGI6bS>HZ
a_)&>PgXe3?\74MJ<+S?D_&?e[5M@5@YMLKZF0AOSV)5G^#.>/53a:(#7QeRGJPB
E9Z\0;<Y.9_efEK@^G20&7L,ZX_8)#Lf#U,9Fa5Jc0QU\M9gYLeQV2/M>1D>ROQc
M.,B=E\,\6[+O58SO^MCSRBNDU+eMU-(.KV6FCg,(d\0M]E\+eXC4RSddC3D&_ER
4DZ85b=).0(QM](\=UL[GRWI8b#O\(<cb,AWJ0B)-Q@]4^WA_A]N.H8f\1Y;cd1J
aN@7cdHKRbP,)O/-(X=(NSKO&SG^Q60db,E=(_eB+(f8-U38=&@5KBT+d-2;=PG[
f0E:PYGACGcOdeFDWM]PZTWAEBb&,EP7<N72.3T\EM,34:FTg-TJYVB-&N3feAM7
OO^B1B=F96]cB&TZC<J[:(1G.=Y.bIB(H\:PRCDf:I#UGU[W+]2FPH93>UWF7HaL
R+F-AEL8W@S><;#ZHW.RA2XQM&)WV^,ITbZPR:Z@PK<GY-=DD2Ga\1GUQD[>M>@T
Nf<<cH-78Wg9NX&N=>^E2EJ908R^#HB\3N=8VO?PG=_Z-_.1/S:=\23J@L?,1KfQ
_,/O]<\1/YT3f^D[D5(.R3&<<DYRIH/+TcJS3LVM<c4NEL8@@#<#C87678+\?9[C
+H:[HT#G[)K,(-F(S?@3#>NIB=F17G^RYUT;(\(UMfX^g=QYd1e/:^^N6E<E\MO\
/EZT\UW,GB.^e6T4&@RIf,A,Ie@e,[[7QGae;6?9>C)0V@01(=;4NPUSc9]OZS9f
8K-X:6;J:aKG^dRBQRW^ba+]I[4DQ2Uf<^S]MgDfO_4;QOgAT#240]X(=_H:B>=M
SQ[N(^CMVGB2S\?5cT=Qf+^bO/g(9c?e,=WS3#e3C7VB76Q7_ae5eL&ZdIOZId22
6&#5K3@G]X_4-)S:bTT0I[)b7[MbeG@FC)#W=T.&fI8I>6BcI[53fG7dg+#DQ2Q0
[OeZb-USdKCdWSD1gLd)BW&TcgE&P(&d69)Z\P]70G5dFSbe+LBKY\G).;FeOO]I
<[W1SU@?[@^BC8@N?T\VU9bgQ0S_O>(Ze>EE+cI=Z77<?P1g&?e#LAX(M?S7KP2O
[;7V,F@fMR;BLCUf862=>cBH;L+Eb8N:_c\(5-NR[J>SQR\M6)SfPL;B.8\eeXVB
,d@M#=2gHF]1e);=Q3O?98:4+P5+\T-==)ZS53/JYJDf=QUbf?T3WVd7:O5U@AX+
2_AC<,df)><2])cQ1_Y\X4,e6Mb[aS>V_QJIJ,bU=))AC)JIQd^69XdQ7L__6^XN
XB8N?7=a&@>BAY28,@CUgRA(64E[A5C/6NZT1Rb/^GAQFf\:CeC8(^[S42>K0>)6
XWF4._;/UKQAc;#J1F([0]S@XNePF_]]-a45XK-.4\5f;Fe?-(2DYS,K,2XQX6aP
/0M=J\]KGQ=0MVTg-.S>=IO\&Y+3,3/YLeB@@7CRQ\1\;H_e;_6(g^#8?67/W9a+
^O(87>Q17#\bRd@C&a8fA8CA.2,TZ8:[#@I0-QZA+7IPb@DU,eHX@B^2NANBe3,K
VQV0]+/&]Fe2_4TDA:3RPNfA@2cg\&W^B[@;YR(g5=^M:aa/Y^.9:Gc_<XbZQg\5
GSWP6C7,TH4H=UK=@\+^+/CXbLb8Z51GUGXd1S_N/cg71NS+gS9NUDf.ef/^Z:[F
IQ+;L4f.<P,gH\6=?32(e>;eV-3MOT8dQQ-ZJP6ecCdg]14g:CD[C\9)3.C,E\SF
Ac7@R0\GD>=A:O:?.O9SDGF^SZXAN@gOfKLB.=aXG)63aOJ.:4R/>M7:_[V6cJHF
QX:DNMIg7>5?7b5_L,[8FU[-0(W<?,NG_YITNgJ[]LK8dMf&ND,/D6OFMc^M&KO5
6M7[;GDXL:V0M5/330BBeSFd0,YUBDE[@?YL-9E6<a@fR0I6<VTPFVF,1<b-^Dd[
]g)ASI:VZ.(2F+cf++5D@_#MP[JF)-BBL)0=I;R,G=We1#3O=BJ1\1eV+3[]&Yc3
]XX6,8[gR&YCDf=93,f8Jg[Q:VcNU1;>05OET+6b2E9W5P(c30)bUTdU,]b6310d
>R=XcccdFbcZIf1+GDE&9MHUA8I^W3=;-,NPWE0PJI2F&9=CLX67-.&S(;>0S2M;
Y,_I)G#e8\E,(ZDcE+;YP)Z6CI,)Q=bICJ6&)_NC\6V.G#TR7,9@&0d[gB,UD<dV
]G+cFI00:d0MQRf/P/Xa-\M?M?bb-MG17Z\VK?^MR1^3DZVHB?ZTGcN1\@GLS.YU
V+&MLcIQ?7SJ#J1W>Y1(JI<QYR-10G9d8GC(M0/V(]U\)\[Z2A9+=#HSO@XVA>,X
EH26A_W<Za7;RB)MPR^fQIQT>13e<<O[M,I[J\T+eEN>+].c7VX67UgYL0PEAK@6
UUSL+=W5bD-SGGW+1IDRdO(/4c_fJC2)E=C#9]0K..C<)ZAdAdP(=]GN&O?BULD@
\c-(c;5EMC=+(AMRYPgZOQ[cLF0c.DDX-R?,HU4SSe22H>LAZ^+FO?<)16GO@(UM
,b0:d_4X+=.4RGY1=CCT[#ITF]H-d0,.LUYGG?K#>(LYK414N+Pa(UA)F>^YZDC_
KY#cK.e4JgQROI]11IFO3d&)e?0QZ+Q;CV)dZ&gSa75#.CB;b0b2Pe[LGK1(I-[c
MJd9C07Wg&09U=;20O(CLJ&7YU(J\aL:=.&aDPEL-M-XRfK&EYXK:8#I;9f1;Lc<
AJ-E3>\),^E=6^d_>10;U48?e0aDY)F(2E-17ER28M65_7dL3R30#86JH=EAUacL
<US1.LI_^Me__F^NdRS8AJ)A\LI5(0-<SPQRJ[3fM>^DY\7[(<Q[HJQBVcVf[F\?
^<CH5BXeGE[d:(ZcEE245F:TSJ->.LH],:V,::(eV1P/T\&HaHe.VQ7G/]BO4#0@
\g0[^6))g#)QdbSXGH6X?,+\HHE2-K-B1-=CKZQX@2b;(Q2O\UB,TB25#&)N<F<5
B^29,D?Oe-?T+(]B=+,7Og4c/8D4>&_?Wf)6f-&Q#DF?.X),Odgb#M&b>4Z9T,YT
N(]+af\B;:KH>(KPMYg;OPY4S^2.&(WQeP=8N],[gD5cKF\WT#)5G0^DFeS:9f/1
>[eNB)<B.#J[1ZU[SJ;0&3AXaX_EK2HW19aH)L1/GdA<CY6)=gN5SeUPE>8K92I^
+H69XY[@9UZV^)dCdLP??^F+?8=M?\E\60LY@M??4+e?R=F6:G[BON4>=1VBc)2P
G^:EAcf5[D=]\d/Q#X;g/1<1>-XKJPV&-7KT#>NBG:N[U\Kc(F/EMaeT)>cI)A7W
/>-,/?CE<,\1]/;TOW6L30DaafD#5P32JDLCNK0?Uf,4NJ]a/[>[KFYY.g.A^7=8
01dQa,/]_b,fKSF1Wad,I-#NcX5Hg[7#,KAS/C:G>U:<^?B;7,E:?ZK/0;KDA2CT
HPYH6WZ=U:]\==8W5)_(Y<8UI:;(Xge&U.g@LO7ZTfcBI2OP^Sa;L.@EU6C]_,NK
?MaGfH6Qb[U[FH7PCe63&6e2&YK+88L.eP;1KVf15\??#PENOIg(e@8>g+-BOFNE
Y&VB_=UJC()OG.4f.4eeLTID5S&M#6I5R(/ca)_OVf2aca)2,#gKc=Pb;I9fAG2+
d6#[W[J(5+d==2(+_JfY@a(T4aaMG7a)^6R=#+fTE<^/3caI.+@=+>Z.b]1^PV9N
/?b+\(=9>N[d906++Z&cfg,\)ZLG[@N^G0:/Hc&)=5</eH]LXVc_KO(9-<@R42JO
E4/ZX]UG,V2#)f>PI_eE05A(4WAY#X^.;77_J_J]]cVX9.D2.ObcY@D)254_@ZM9
[I6YF5DX3=f=M#C5cE6fS0Vc5PWA>J?^DEcX-g_X-eKBA5\cKc;:^?LQ<Ag0WVJ[
E;#>+_F0>TAO-bTCedc:><&_&AY79Kf_bJ#^N^6+1,@Z__46W_@a(?Qg;GPO2XY\
X,=eO?)B&.95cK^RTc<D4dSA]=;Jcg/BdHHD<T5NF.LL7#Q&R9SBTZ7DCJW6U,D,
QNO3a.8WY(9-GBJ0R>#9@L?+.>FGQ;AX;P+@N5I4b.8XKGeU07\gH>R,T_c&,MU5
ZC5TRZ=-0f(GHbIS73)Ze>b0EBGW4^.<KKRe0#><=]d0:63.H&AWFH.F31X\.ZK>
_7FV(76^2[JD8;UL2EXY+8PBcbNWW.?RdLS;GWH>.LgD@3>c\K71gSg7E@#4O?Z<
\5#cg@77S+/R:W\RF&LB@=bBXWY32:5]bONOdX.Y8#&+],4X[QUX.<N>9RFc0f78
O3G1CVWeJ4Ue#@/C9FG?TA0DL.-P0?F6eT5CE\be0EX\U.<VN82@UZ/[@:GDO\fQ
6[?_2Y/S,EWb4Z5JM+aTYW7/e+Y[2@X32>BPHJJL0=B>14Qc7Da)69[=F(G/d803
ARLa/W4OHR80[S168RWROY/5977]\-B:<\Z.BaR<V?L,e>eQ5XSR:B/(9_4[>O0F
S@1OW;JEZW]P_U-MFf\R+Q6&\_83B&061AD_QSSV.4NSF\;7FTYRHY63#K#:gf_R
0,+6<S@FK^4-d_gTec8d46^(U=^aBJe.,QDEC\/)KeH)HL?-]/bCTU>IQ.T#AOEe
(_?V#[/SZ/MY(0)F6Uec;D80;K\>U;-SE-<[))82]XfTOfY<R@-8H31QJPIS=Fb9
eIL05D[][#]-:F\Ic@QF^#8=N8M&G1]?B?C+AfT68@f[(WD^419Xb5MfV?3P<e1F
O&,@=X@-bIY>IJ\a8U\UZ&H?K#XQ=&g_KC@b6,05@)GMO.,O:ZY<ZT-@Y3P0?f@_
(97e#Gd4@KPb_eIC:DXIO[UA+W4UJK]P,8eZeR,7R\)OF[VHC:.F,Z23Kfa?Z^HC
9K:;MX+=]Cf0OG1E4X@Be-U4RJ91;-OJfJ(SFP=Q-=BCS,A3#6]/\\3&Lbe[fML5
HcN#NgHMdUb-([4-b9f^&Sfgae=6&[ZY;J<&>NDS:2,=;];e8.\WNE4I_^L_DOe\
X9E4ee/,I8F&HI?Sc);Ad@b0Y=OCKGOJYU-eJ[(J&@e20U1?5G\3DEJ8;>b\N?35
J?MD>3?9YN-SJITOW9PD.H0,ecbIKPXPHAT@(Z+SR3<P><b36[K;@^:A3LOG)b&C
^(^Pg&BWKUE\e49SQ=JXAO.A82;7g3e]_?N(BWF1A^P#T;:aIU6HPZ-#/a[VY)VN
0eF6UAE2aed\X/\2fC6RP8TV4UG:_JHMGO:DaNc6b;R,+CP&gd(1KPL.5]?FH9@P
4<:9@U(6-LW7.bQ=RJ3Q=HU/eLZK-Ua4:8bB=GMgg40Z95M(.[DSFd<bGGA8F8VQ
b]GMd_^XRP?P<[I8[JAH&G6Z?JeU<8NZ5<YTNd(A,g4:,(0N,P2D4G/QdVH\FIIV
QFLcRC&O,0I9dNgA_WWX#5YL:\d>aR--L<S++J;V[&(>6JF5g9eK5ZJY#1W@F<#Q
LOZE]2ON:3d-0JW2MJU3JAI>DIOd4RX+G0&H(N,]7X@NQgW:LA]ea^M<B.O/WN)W
E<[0#UQ,M1=#BE_CCNU#a5g;/I/<L6G#<gTYWNVMU-V+eDBQb_)#@JS69LCO_WXY
&&dg-PQ6F-ZK3J+Qc/9OST>P\.c?-S+5?470cQ_f]c9T9IBJ:41GM1HM6d]?#@X+
c=@VFdS&Ka8f?We0C?FP^TVZ?\7GUB<R<\L1W2,HBaT)R01P-HCc-JZ)T>(1bD@W
KY7D(NAgMe+bT)Y;dc&70/QbC2QHXgN9aRGC/GQS,K8G4=?ZPG^;8:?;Z4\ZNPOa
>V6^fNXaI&_U=T5f11cHM06)/PF;]AX3W)W=bX7(XY.-KR[=#19a8SR:]3d[7S<C
X[NU#1>..0)Y5UM/T]7NCIDcDN_9B>>.VZ2M&&KEgXc75dQR9/#A[0@/<Rf)F^^\
0-X6RVOf#>cJ?F_[fK3-CD_\6^cXacYJB<Je1AO0\F18PcgN\d,Y/[8F[DX>QGD<
IX)CLEgUDM(M>9JJ/f/gPLb\/]9aHdD<5M):+6dY,,a3X9_AJS^CZLd37W?bLNd.
X9@92_USH(QB5^L=0<([P5Hee&T@.DU4#7P6QGP2<?MV&[/.2V8BSX(U08VDaS76
)Y#WXDI^d/JdcbSQb#TP.^SFZ[O_2IP_.4I4S07[B:gF5@&e(^9Q)N\NG/0ONc\C
ST@&LPUPZd8[J@V1R3VdJ0;^-9H87BAGEZ38F(G6&8U)W>(P\F9aM\<V^0Kd[1C,
7#RR6^eIV@UT]1aL6=F6R81,HcT#.Y])7@]fTSWaME4C4#S&4.PA:VDPLe\RIE51
c136Q#NJZfCcQ#O-Vb0RZ</:>G-K,(9d#8Nd/d,cULJe8<?X-2UBCc<1D+T?QFPW
\X^Z(FAJ+SPGdANM=C=TCXP@d-\aYW@_Y9YJA&N5A2;_06?(R[]>OP0F&c[=cVgW
JP/_X0X#eGGC:;_1G.4,bd-dZ&K?dQ[4I?WZFA5[O3Z>(4M/S)N.>gaT0X3.>5KW
2?F6B:1VMO#OC]-C,?QbQ/W?-JW>>5+9C3XgT1S:\/7a/OfaA5G81I)FXPceGF.5
K:)a7I\gL)C.W4CGbIK;a9BO&/3JJE7AK&ZD.BO.UeK,:0D.HEfU>[Y+DKRQ;e0>
ZR(2A6/FFFb:Y4R(e)U^J):=d&4?=[TDYO6.IeaF\M=T0g2PeSR(52B1:GfM;6;b
fN2cMd>=gJ_<S+6@#UWeO0SYTPJ;SUHV)RBYUefeYaG-91=2e=bWGaEDK_dX01]W
H\c)36Dg]30QBSZB9X-J+\@\e+;bdVQHQ?B@/-2\R_SL&QTcF@2e?F+H;HCI)\e.
?_YPbK\CMA0GJ\8>25#^(IS1bRY@Q&ed8_b]\a0.@AF&-#2?4R=fFBPB?c.d4V(7
NP+\9I]/5?S@c2YT[XWbER:>e#8a?:FV(M\+6\3,GNZG12T0H>GefB-^Q\b39]/O
[R-QeB7bM<cF(LP:4M6#TKQRZfDX;LK-R[-E0S/+5N#9bS<+JGbR12K.2YXB@8_A
4@2^U?9Q^4H4H&F[[7fXUDZ5]eI/<f,ZDSY5K@d_XJ=D?4B@1Sg#=@aVW[=b^RN,
dEIccB3_Q6JZHD#?2O;ecYK-G^6=\>:O^ELK#F6Z8&S601.WYL_W,\1a93+9g:7,
=]V4_g4EN_[cB-aG,.,-<b)+NIA5MLVf5?;[#;-V6,>><Y\dTCHA1-;,UT?0#1YC
AB\?\5,N#9c7)b>:2)^+P&MG5_(?Me/QVa#VB[5Lb=5.7_5feTR[7:M+XMAP9FZ?
c264GZTB=56c72NBgP(\IU_gP)[]0[^,L83gSY&g#AJ4J=#.Ef<P^R&JDeW<MPfC
4+M29P,[YH6L&CW6gX?6AZXOE<a2B<J2@JR1S;OKH9#OWgPCbabBOag/<OdS>a)F
U<6g]XILL9@fME\DB,(P3[=J0]6FAfL?eed&M\8gCUd]WT=7[962^;8-NN-2LRbY
)EST?e2&<G9N&7=XcOY-L#L#QL<5O7cB7K)-U<N=QM-aM@+Dc([4<V3aDg92HQXf
A\f(0g.<ELF.[d6GF67Ab(L#+^7<IdC?Y-aAgaX&AJN4&,gLJ0D]1KX<.g<8/1c.
H,<KRJ6_#CH@cD&X,EUR>>OdFg(RT4FP^BKPHc(OV-QLGcBH&@f=JBMfL87gD9L6
4ISRR0MW6M\#(5TTQV0_+Ad9W<S#C8G1[18;_Te\;bXe892_ZHPG+c)/1HL,K.9N
FK>\AO\M:-32HGCf+V>I(c+eSN9W.F\8L(0-.MM(JO,Be(K#0@-aP7CP1W,<E@I2
_HegET&91TE9YMQ?&NC9FTY)FO9,=WQR(LBdDV1RZUE8D1C?+_00:c8>^(.,D<XT
7b]d5+SJ3M-9H>ZfLdUPLV<9PZ\(;d_<fJC;K3-PN/:<aH:b\FOV<:de(NF<G,T4
T]&8#aJBB<UT[ff20Q85AE88K:0e<23YAdbZFCOX;OCM)]WR2>W[#-cWJ]P8ZG;G
\K;E1>UM(@A0GM_dLL(E]XNATX;P<CddCfcaD,3F0WL6)YB^#48NX^eV<c5Y<+Y=
][.aC4\C,Ag+Wd6J80gBa4;@]BLPc^cd#ZIBY,K,1VNU)2CH&I@XW8=^H4/C1Ka7
P322RKNEbCUMI5.#IA@7/fR]Pg66M]gI/SA_Y^(0M_R-H3OOS-.UK=BfS@[5T=XZ
g,<RHN#)0C0/?X&DIIYdY(=HK=YdgF,6aJ(=4a;0>^]VfA1f>Z+H4IJ;]05ZIVWE
.G<IKJ.X/L<8IE^T/CGC\cgdRQdVWY43,P[C0YMeUBEf]+CFRG,^BQ.CC@P\.\JL
(+BCS>e0\MIcW8I9(dOVTQW>7K04LJ:/6c^RQScf#;T1gKUHP#d1_F5@d_UL_@]R
?>@Ee.>4/9M2QIBcObR?<E:L;H8DZ:,F/[<OCdN\_G_;?+NO.&T8dbLFD3O0&]Id
<c\NNB+Rcf@=a4@f(2d^4Dg193B-I1JS/(3U+UDcX6TD_6dae)FO>e<B-8U=#7>Y
AREa^?F8d4F/&>e?_]E#MeWCcW[KcYD-\^gW>Na#QHE@Z4La<#Q,Q\>04N[TTB-G
J:+D5(05)W:+bV#<Q3DQ6Z)XBf8+;bfTb=K31L?a:BJYQF-KJD;DM-Z:)UW4ZWM+
S_)9=a+07WMEdB/?G)[bK\^L]X/1QAE(8Qdb\.gB5(JV?:#8f)]:P3^DDZb@?G>H
/6fAOB334_Dd2GF,I_d)8G3GGBd78JaHX\a5B>4GAR.E371bU(cQ?b7+KL[:UBf,
.9\CVSHCVNE;8Z/JP;53BZ.RYGB6GGaU=4>7-^e>#7JGSB<Q_^Y&<f9J[A;\XW;C
#.<(=8d#=&3V[1@b2cVK#X-RBd.,1=A32(]+5>^KE0[EOG-K]Z\A0P5M([OT0Tb^
65e@KDf?F\Ae5XfU]8LUIN;]cN/(\0/C^)aP/3HdF-GS7LFG.-K:G\WgAg29PWP_
N:e&aAaH]LeKOM?<>W?2UeT7@@-[H@A#B,YVAQKPVI:AP#WP0VgPKI[)]g\):3XV
/-#Vf0N?ZD=:MPU(eRQag>9XU)F#<Z@1=X3d1WC+4fP1-VGg^f:L6YZ@RPJVfWY3
^-8DV#;N9:L@cOB&H[V4U24B6e3<(#NbZ?c_&f884W9?L[Y2U&=<a(.GIYC=[>K_
PD1XAT(_cW-U5)0-OUD::(F+KJ9S,9_&3WbdMUUP\aMKAaeAW684LZ&WMJA_=P.:
19M2\.Q^\2PB1UdMAc>8A3OPXW]YTPV(DLXU>g&W?M?ZJdeeE8b0BE<K3ZJ+N1(c
1S6NMXXQ-GcO6O&17eKU^]_B;^?\MOA1,7>2R\41PBfQ<YcbdZ1I3<AQU\D<^3e&
O?&AP).\QP?ZIDCBcEQ[MH-[#Y(J/M_KBR6?VJ-XX^Y+X?+;]&Bc6_C[Vd,\-08K
U/4;THRe>XC#bbY(3)eVD;>&E+P:DM)-)YWg22G,2(OMWdEBS9P.X:2GD_W8@]gG
E/0C?:-15?T@.EJ;28&IL.2BEa8OPTP+/BPJ=00f/W#HEL<&f/VScGR47>gc_E,<
25R)WFSVVe9\<+SHX+Ld)2UCK8Ka(=AHEfI,?^ZX(F8[)10Gg]J;@K?d09aXHbcY
@YM(;?X[57)0WSS7GR7VF+13:?TZ&g]WR^_3A)YNDH=fC\L[F:F3bc;Xc/f1^+:=
NBfI63>B<TK#0;dB30_TXWV+-7/U&V0;OYO:R>R.F^197BeCa-8\.MQD.;67G:4>
J1279J-.SFN95@0NL/&gJZMc2N]M@RRSJ-_8=gC7F+<-7OCc8dTL-2GL>G8BG(<;
?QVQ7WG1&M2g70#EYKX@QF0B+H?@IUDN+M]c.A-B2H[Fd&YVfDd5>+cR:e_21I2-
&V]^fQ;eY58>d9UD#GJdY5#afaEf=FAcM]>d.YX,)7+L=Q[b#&eAaL.],e^::9_Z
[VBF@0)2fU8RcC3a:EV?LU8652OG5\1G3IXdb=<&3<(+<4\.,>_7MA:4/GGG=@=#
a6RK<&Vgc7WVONGGK0d2D_CS_X4_)I><-<CZF/#HCDJO5>JE+5)4@^R^EN9a9DTZ
]1TS-VbNXF8KgD(-0f9QW<,&b(CAU@=X<(:->US3N@LFL,SLM7D2?P:c_O#/^0NF
T&GFfLbW(2T@c(eO#<Y;b&;@??AIBP,VWX]e+fD]A5V5fg<<#fg[a:)M3)aNEBf]
G>:ND>J8T#XN6^1_(,17S^1fH^+21Gfe;TJC8;XNX=7#RIWUZ5fYO&TaZ6,42)dL
LR:Gb=Z/Gb8++KNKBW,SP^[QH[9aI=WKZ1U=]+W7,-L_.gYb3._@CG&O2[GF_L>V
]/P=K?9UW^#ARYX,RVY:f[PZe)UVIc-;XgU@:48K_ePg3?KbDN_7TT#I(6E6A=G:
(WYH.,,^0O0fa+Y+A>34:1)&UH1>8fOT(^AKCA/FD\DTA\F[1d\SKPR5[FAe>:2)
?>70P=HC?UA<VIL5V_Q53HRQPD?^QHF5LCIeSZ0d74PPX_3;Yg=1NHUNLU<)eM99
/:@Y[THJd;9<D6G7DAR-9C_/3)@/(XYLO;;_?I5,Q#1f]I&8<Md:GdO>@-QfK:c&
66N11J(BK-:c4.]e;&55;#Y^#\NF@4LIeCOB3Q+H9bgHN..af&IGE=e4?631ec;2
b0]C&c/>.6EP@O:TE:T(_C5AF3/V<(e0]42H4FV;KCP4\6I-M+T-U3/VI_L/J;/5
C4+Wae]T[Vd(BOE[aYg\5ST^f@BWPI5ZQaUTSHHV\QRU>FGX(W4;YdOfG+LMb<#>
YO,T(B-<X<NDA;[M,+=CfEK=MGRAa29^gf(2L#USd(?A>N<=R\[.LU#TVCJTg,Gd
=M(N(?VgS=?#OBZ<?SCH:d1N&E<,Za?fcUJaD6Xa32V)e3P^;?.N=@C06gea.10I
XB:1-:L@#>4.FGG7N9B,TP#07C,eATfHY5;cQLC)<P+_)=[e]X>?YD;9[V]HT;-#
4P2F0<#I&C#;4WBW81=O.ENPQ1eE\(,?@gSg=<a\IC<bTfDLDC5NUIKXQJQI;0BE
;.)Zc8#+V5#;K9X,YX#/<\U,?)7/+BJ7cFWT>E,X]1T/1[f--a1#6S0>9W\e0A[@
QFL(L22WTUJZK0RF4&;cAJI-[Jb6I;S35[I-;IDH3\EWNbR95?\ZL1?cLa+OdHYY
HQ\]J;00J#)WP\YQO:>?VJ0J9RDY220#V5>fGgC&DK,VD]#dA=+):YSUdf(2UTa:
A&W18Y\?S)[7P;Y#X^Qa+[-=cdDQL_+@dWND.&&\W\OX@RS9W3]g7a)&FP.b==BP
@#6DR&6UB^8La5c-+-b/F,11@7ZN0[^T+X)>UXJ97JYEdXRTFBR>Z[<IUMC#M(8#
>7=6L4?2\Dbb2N<&9c^;]O5^KU]F95PF8@^OMZ[+^L6QbVO#:1IaLW:,35N[ESKM
aA)e;WDW<4Z>JT>+RZ(C(_G@DE^MBdLPME\O(#:M+-+g?S;8Y12e>S2M_(JEWeKX
[.C_,JF5BM@PZ4WcW3^We?N5^1>R@e#(:Pa88H>=M;(#Y:&Oa5\PfMMMS;19@dVb
^G\,de1b2d5^[NKIP[Xd:Z>?8.2^8\YD[O7ZVY0:&21(QV<HQbMV]UBdWbd[>)7g
1AM--Ab&RQ_@1:FYfPM+<DMEda1b7NgM@gO?Z5?2ZeLW\V7:FP&I#EN#Gb=HJUVe
?M?,?&I+cSFIGGXQSSB2D]SKK/VZUZO-?.;DUaB:.Y]bRNN)GSL-YJA4(^+IEe24
=_UQJ(dgaW;Ud;R?^V[/9PH>feMK927^RD]41AOEL:5W.OBfH=-b<)GaEVWA;bRO
fP6.d#?<JFLRX1Je.>_>KU&b=V;X5=EAC::SXD+a4Q/,_C9YF@=MSMYX92R?&eD5
/7V]E.G\S&a>EIMS6#9W1X8^AHT)PSb\8:f;(E6AABNEECG&,6YX[ZcF^ag0SV9=
9Q&-J+UD1==FU.BI;E\;2X]3\7]P@a:cQ28B6;&H)#F;]A<f)c=L6K2f:Xe)1YQ&
.c[B,)6YEI)VVBZ(,<.aOKR1Cfc+GKU]&4VcXDYN8>(E:HNNK>>[NJ_RTH#\CO.Q
C#>1N11GHg)SKYV;]NF2Cf&5NIM_A20XG;ScU=V5NJ9+D>H]AZ=,MW7bfX?NOYQQ
J+]A9G942Q-)gGQVS\+0+MJ(72\3U.)<@@HNFT^6d3;HT[PJ:QDAJ;+Ka3c9V\<3
JNON;a0S,.f#c34e60>0;B-AOH5,T2M[H@e6b3BAA:SfQ4fRQIPT^/4?/Y:M[^dC
UfC<2-Y_f]/(SX-Z#:YSfVPGFPV2W4,,EJUd)QUNN&6QQ[]BQc1WfTSK8RH0C6@5
EG/27<@V9=/E46Y@)];eNS82J?eg[Ng0<YLgU>K:X+^CFFQbARcg,e0.]-0U:^b7
?OXKK;\FPKA.g4f4W-N?.+F&:;9M/[_4+0fLG^PZ^0ICc6#WgNQIRG_a2XCEaBIf
G,c(0B]Cfa7MK__Gg+QRL]/78,W(N(\?Afb2MgXQWOJ.Ge25.E5N-_<[=8a,I)P(
)@Q_<5TSNgR:+e+eDHBLXT6TK1a<HUI[12E8JRU57aXSEQ9=#H\D<?5/1HML3cTV
\e)/(@/6>7:eB#VAVCBT?@gR5.UHgJc@UC9[J3;.#-+X-d?KA/>_<Wg8S>U<G.DU
JXCS3T\&,/&,6(<3B3Q>,c)[D:P,^7>gB:5BALWB#F-W0D.Qf15M-QBWOMVFg;^0
bH1c8E22U(A)2WeITTbYb=A,)XfJCB:^TD-EH&?_S))7\PLA?@T#0^f2R<V(ZY-1
QQO.^(1eb>2/P25,Y@:J_Y#]GcZNRWOHER-HW7EcQBIeWd:8+8[:TM2aUA)2Vb2.
9d-X/HCUb.40+eKGH./VQM?,F7[E0R)N9OaWJG2Y2.e&L517e]]_H\XNd^>e6^W#
=:>AE4H31bM2XX?A_AQ;FB]3V\NQGX?1GYR[\97FDLF.RB><.HBG3)YQ?QV\&#cM
VMdfC>HIN7C8aILe;V-5-f4ITNENL;Jb\JTOK36LQgSYP7-.,UIBbR5J?E]g^H,[
9;O&XE].PUNB.(_TBfCP<(6F=XY:6eWc9(+_VR\19O+E]5b#P<Sf)\ag(JTQT;T+
-ON.BYGSa\M^c&K[9fLdF^M^b(1JJE2-E2_&.]=FB>)RM[QYG?+F9DX1FL@G:K@K
&5d42E])c9+>5FM=G9@US()),=\]bNZ-H=<?5QLGcTY=aA\/?I>aRb>:\NCaI0d7
YCVJ248e1gc<=A9443B@=EKX5LL^_1WXUGSUYL8a)UKMO##OXZYbHS2O<44)bOXE
Q2eYc\E^7D2(AY.O,EL,g](H(W(a>F;JJ:)B/D)<SOH3;J=aP3XOA@;deA(C,<>Q
<DEG+&6@)@8)A=d&K:L]H9E:^f\:O/5e8W=&dFP2EWb/f9EbC;LV\<>1K[-^^0;7
^<UHVdORJ8Id.#bTH&<4O_fXSRM+],91aQNIG9)S>P<0\D@a9?D2J#QB&9Mc/Kf1
<W_MD;_9g.J_N3[c(5P>1&MXR#)@/M+MB-A7.JO,NJOHFa6^B.0&T:WMMZAR7beF
-MI1.GY8U#+A(f?UT0KM>-HQ@dN[2>-JK8J<b)]/=GfSd76#-KI1;_,QcD((G/3;
<IW\9aZI05_U8UQ;/fdb<^2V<.M)ZP)VB62bf9S\@/_O0E8^dU1J>LeWbQ1?+FaR
dXbODcABC4?8L]T)U7e[VbOf7=ZYU+03Z&R#FGSCf\DN\(]EOf4V,9I3<=X&5RaB
=4M6->FQ[;QfX76<P,Z409L=9D8Lf\c26_D8PcG<WEQP,4J.Y]ZcEE]SK@@GNX>W
F-EM>)d_3@[d/>64A<WcZdC_:\;d<)X>E\Lc?PHK-XX9F+T9\AgXG3K:^]+.L68^
;8\5M.]YQO]P)9XA0<G;YXY6:P9UPgUS->FAESbK_YZ+?)).9Z)Z=He]F](HeXQP
Cc/GfN1,XB6H\]@M,#IJBWV?1([R);:bJ05C,8dU(8/BD2GB<ED32eB(;,?B3aK1
ZcE+,)(4:6SadFB,]3)\eG3EADZfeC1FKgS@S_]VC1>AaIV+GXD((?^K@cI\Bf@A
A&.Q#c=9D_X[O#X/P-Ea@eNe0LFHDfX]E\Eba-J)QSCOCY^g?1?RBW,W0^Ab_5?&
]3VYQ:;XEV<LX=,8e.f,[=XB0eS)Ja;0;X6dTdU_Xc.ST(DSGO?]]-DG(XD9T4?J
PQa\WDe7FX^A:>c\_4S)\G1Ma\#@.:\IF\3E-Qf[NLSF7]LEO(3[2[dN97+BE->X
-T3>0:M/S=dObB1X_[T8MOVW/(CWRS.1+N5CW_bT9KSO>@>+:X^RRD+OG\=/LC9-
KdVWbCfO8Vb<WUU5\3^4G<0DP?Y<D#+LN1>,.&96BHYQ_S._G@WOfK?U2PV0]O=X
b99]2fM&8+<M41Qc207]07,T?<M7W.D0L?LQ=8^GE8F9G5Fg0\SBZd94+N:(3N:9
N[1<cf05>dgbJWSP#DD-F@NV2#S2J&AfD/\FI;FU\@C:O,6+JNB<RdYJf7<cQeC9
(#MAR7ZA?<Ma:&>Ee_)\KMC+.DN[9ULNT[5YGeE_W6ba4QAVa#:g0YTMQ+)A+CQF
OK_9]gI3K3OFZfDQ+Wfc]?X@&/&a[LP>A5LLGF9E7<K;S2_L8:77T&H;)_9Z0\eb
:]W8]:KGHN\:f\]N@-g<]DaDe.=L=,g4&O-E1d3T5faG<2c-NIU#&B2d]Pc0\F^U
aa\SAMASDVITD>T=0V?(JB:#4a:YV+dS&NRH.Ld=75Tg54F&eI9Hed9#UO>-dBL:
KMdXKaf]&f/8>.)b?-G\,M)b-\#ATfc43JY+,@=#QM-/cbMdeQ3fG@7AP/7f6;/f
)G3]S,]b3Ee<<ZSefB^A8R(81U_0FgJ;P,5]YaPgD=9L=#^<]GIH5B&<AL8JTgPV
Q6Hd_gaX]YPEK7c3;>7Q;TSP\SX9I3CM;K4@KKA_/^,AR&RZd?B/:03>]gTXS8HL
;03(60<AfaHe@OD[/95VJ+K4T^?[0[Y<R)KN5CcDYT\aK?9(#2LH1Z&DF]P]bSD0
Z=>bLF/+AZ_:4MSZ6=QD[gG5CY3_\+QMe,g+9O_,S-)]/D^SC[#eNVC1MNfJCf[Y
.?<U^BM=SQA@7=J_+].Y=gB_g[(GB>ADEVI;H(>f-+;CQR6(Z8@FVT)BAL@#X(\L
^/8CJ5f;_S3-V[]W].P[fR2??Z]&T9R6Kc5004gUaSUF-LFNDK+Cdg,L\XCd5BKc
0_^(db1KV&3.0?1[JR[A>=@PO8PVDf@fJ7cC@5MR&Db5Z#[Q6\QeFKU21BJeE]^.
#>DT7TD^013U3EW,1<]Ye=71RR)WRSUTdYRf8=V+,_Z2UD:\WGB5UG3eDDH=.WaX
cL30WLW[=WaGEXB5_CZW0<>]LeRBR#[M8][H([@-@S=:DI3E;8fQ&T=;.=2-8;1G
+71Hc:67]=@RC[>^:X7^+1JSXd4M6NV.8II7)\HdGV-R&.2HM]&cdFP,d6SF>#60
1XTB2WO?c?M(4^+0?+QOL_cFY4AEP-+JYf#H;BA?,UK9ZJcM232IfgHR>TF^A1/L
950_50dVg.<]Fg>?\0WTbG\/d[YP/7T.&7:gX7&L@,Y0LB12\UTNGPeJKL&H/),@
Y(1[[H5[8E/F7(NY,JA9P6Rb1XC1V+XUO:f,UFe+80#]<<_HU0JT<SA^--K22[SH
-,>)YU4L=?dF\BTU-SH&PUG0L/B_C:1PaL.WHN6,XL.JAW=>CLgNVM\WIPT49]9(
-SFPcJ)\XOWF+Oab(;XL(f1+9[WN,OMdQ<<,9DHZ:Q3?6A>P))E\[QA,9@.55PGW
1WK;Xg2B=P^C^@0<U-WA;[G>FH[E,.I)BBK#Sg8c;22[NQb4:7Yf@1F<>\.4W8)M
<_A]9G&=Ca_@F7I:AA5V6>.GJ.OB?&.b#&#Xec45OG>F#dbe3I;LC#__RSE,+A2Z
Y<\MeE]8e<dCYX0DO,5gCTSP@):b4MeC^eTBc_L.1@&_(Z@9K@0X)7Z/T\CF?4UW
1ePE)E]N0<TEUSRV?WOHLQ3#QJ(9JWa3L0@:WcTJF0E9d:bEQPT;<,6@936LJN;I
;_ZVg,\_PSU.f(5H)?e/C/8XP77\A33^dS#@6_S\LE3O;FD0\K7Q\S\:PX=dX4Z#
RCJYK:)Dd#O@L@T8JG2X3RRb-XN-.W0UZ41E_XE?8:cHG@C,ZdQbTXQYB\d15e^(
AB(TB24<D:]>S5STVLc,bN@J07X(S,K\&8#.Va/_b/)TJc-?TG^I=L2>[IK0W82/
XgIMN&FL:P=;[E(^CI@8ZPcVSSTHT#(S4C&a3R9#IP;=dK?P9RQ8Q9[M<=3+8fZ:
.Jc(f+a-_X?&e4_JH^2Kf<Qe<8E)A#CCYSQE\&I(#D>Y0F+A#S>&TBN)&^^;6DG4
]&H.^#:4H-I:BP09=WM:J+R#&NOKA86--7PV)W+P_K=L#MNRN1g35_Ve?(C8:M&2
8P./KSe2?1Oc^de6-TS,S)/6.LDFUM&;<b@Y:L2D))MZ2bH<FUK.[ZQ3fI[d?.Sf
6;K(Cd?1g><M-KcAAG(f+Eea..#/U>Z7^]&86=_DA(J+UdC:GK\6D<&#+&?^TOI.
(>V<,#5H_(6,S0OOC>eOVD+g5@]0XO0+a82M.JFCC0V1La/(VWb(A>__B;AL&K&0
#fK\3JZ]0C_0]##Y5-dRfM;.FWGC.F=>C+Gd>fL63/+3M>[)FS,/UOW7SgUED7_0
g)cLD2T;\fX^WQa(38\\O8&25XLRZ/QKF#/7B/P>c&/2+[</F0G08))[UKc:>NJa
#.6cIT)X5E6V4CH,5R6AP-NK+<I3MSQS<Se?#DGC/KK9(BEZIT41e-835O44S1@N
;,b:dYU@=)RLSA>eNe^X5@ZKe0dV;Q6#<6T;)V(QLc8<NV@:L.43)/83HM&38>GA
[6acL#N=.KgXf_OH6cL[,A<VB6G]+OZ^252&/d@ZBWH8@L?WVUPY1P>MAX<UTaE0
6RA\dMN69./J:V3PQL1)-PYS/[LA;BP_5>5)CL_80Y2b^a?T^P5fF)ZbDaNR-2Zb
J=;Me<+V6bF\=fA;0bI3:MAY>#C_8:9e1RBZ^c-9\8>Z2LVAg3d)-aX>1.\MU-[L
WULgVa)\@<C52YL[O=[UDbP^BV,6(@-#T<Z->28)G_B#=<?Ka)>8:?a\1=3/_:Y.
V+R,;0NHY0,B0_+KKULJJ4Uf\NSOI9QZ9@:Zf&=7Y?6b4W7A:T5U-L27:/D0SA3f
eC^-Z_9<SS99K;&PK8QEgBEfG:]_Zc&\73F1b?cCZeA-ZCF#gTI)Z=a+N=RZ-LO7
cWYNHUc4e\\&#G<SNEF(?1LN6AfLJFQEV]]7ZEGU=8RgUgG@d/AI(6V,HVTa/UJM
eQY+D2B.VF@0aJ?2/J[V?AXO#>Y0S1V-IZ(H+),HW22C@@cE)Z5CT4DWSb[@:^?T
XO)F30_?CG^?I\V?S5GCFO3&0;I&Z@Qb96W#M9)(eJ4[Re#T(,aI-dWAVGAU]]4F
UV]dOJ7E?@^3L])T(523Ge6-\,#Q;#/AaSH_S-8:D?>d#VVgfdK4PXO5@N&6><;<
)fa<+:a1FSfe),Y\=+(]U8dN,UBcX63DCT7bMBP4YO:gW)<dPSDRUW+Va+@@_4(b
W+9]>.7:#6EU,I=?Y-EEZ+UGB1e=eR<)ggg8O&e?YBH5cQA;Z_[T<C)dLaH#-e?)
>SP7#I)3cXfY29M=.166U@^KF[737S2AAY=@7.c)8S)2-HHL&==360EZF;RC8[U#
3978cL::1XG/M,7P0BdZ@IW8Xc\^cM-U;b6@MY>74d_(#c:_;[D[=O.-QMK8IF&W
3:Uf84PRP>E]aN1=MXD/X#g?SN\QgBIbN=g8MZS9?D)D]H6OgE7@/Q[2FY]9?\86
f74BTMR30;7Ef@Q(Sa.UR_])K]_D_G)BL03M1A29@:2H4HZ)0QX.[M4a^KWV(ZeW
>3V747C6N#UEDJIQ)O#PTGW]KTUEGO43O_ed?<1\LP^_TN25A42([JO,NEf&#O_<
<+c2BP@W(6-D0^)WC4DIc]RNdB(DG:CT(gdTYKRJ<\5_F5BdeA\be.;)5G?]K,0P
(;,[_^@3IB?:U2\IZQUNCW.==G<c\#[->]#W015[RgCKX^^BH@T<YX-8R[^118>,
M@A>+7#_S>XSFV)>MbFW8g6aMIG]0W41eA.&UJX./.NT^YQ_:T>L4XIbP^(T6QBL
;<0ROH?YbV,eMfVGM?I31FE1Z(M=-)8E)^UCa&dd75R01P3^K1X:QS5PdPD_^XeL
7fQW^@?F^<ZOI5M,(1=T9#ZYaXf_3,QBUVG,GH0T.gJ^&L/2;NT,#aV_-O+e>GaE
=g0JcYWd,&Ff.2H0LSd4>ed8)6b>CGUY-+^Ef[SXWH?S)W7.K73^)_;WAZIBBLTJ
=(.N;bZA3@^ADg&V.(F(^BN,cI.[.&+W\ERUY?.AgK;Td,c\,MIHd0P:P])g>231
CL\K>]NMQb1g\UdV;=CM6e<;7#aKUdY#fWf>,S9HeJDJY&fX]/5_M;BQ[P[>P7:2
\(8_3K;&0Y,ed@,0/g5V-R+?PGJ#3G<Y6;UH9--B>:3DP3X8dGOGHE[ZF9MB(HdX
,[aU&3/M7TWa-)@&O@]--G/>M.?Xb?1eUT3c\)0L.7^WI=67]LX#P^X-U.H5TNO-
83:8I(BQ06gQ9>[\D5D)dee=G;aO7Ya7LF55H]?4LVeER/A^0L,1+Ofe-O+24O6;
T-RODGP&E,Z>9J>EHJ@08[CS]O[1&;2D)U@9^gS>_(2#(EA+XM-3AF,BHZ/V#IRg
K2N0XfHH6RZJg,Bg>Q_Y30P&TIb@IE[0;QCB0>-U\AfNRcS&T12F,PaW_-0I@GOb
1&cR.W:;V61aP:aNBL:Y9O7GOJX3IG[KF(CTX\WbI^8@Vfd/2:?AV2RgNXfW.)9a
>T6@U\HT?.S@=&Y2Ga>#Q._[C#d-9VD^,(fO[=Y=L8;U^2^FS_+3R5C0c8GQ0JKQ
AYI;^]AW<T\6J4=(N4e[2Fb+IdV__-N)&f-g7B[dKEQ96f3QA#2V,G;2_@YJX6WS
XJ3&R+65OR9H:4;QN&:b_MS>dA?A1?bX-Y,#C9CF=K@5_G&dU?b=BMK?3<YA_S-L
#e-].N.UgF^42Y)0MZI^,/.,/?7T;gC\<aZ)&Fd8BZNW]8>^;EbO/:?QI)H\;aQe
+IPCG[8Mg<+PYU3(bOfK&M1=4(D)9Nc_C\JdH2Y)5&QZ&X:L5Ja_]CKZ7O^[XDS?
:\ebK6^K\+BQYA(D,#e;.=.,I.,IYI5(8B;7C2ZY#@fL9<:;K;EfYeD(5VJ=QZ][
-d--0U8-S)J(7dYL<Ad5Y;HfQaS(Bbg,--\TZMDDW6_@+1?\.-:#]@I53_D2_=)L
J29\bHIYZ02>YMEKV<)OEbQ0B\Bf+I717QV1BA>cc&OX.e.L0+L=FHZPQC&NK8SW
.&F_B^^MBQ]<e^d(:+NOZaVN5062f(B59aW-MS#CY[ZTb3+9:+-.2T+;8I3\EWLR
/P=fTg]VXJM9-G(cI4ZX>Y;&0O6WD^],SRJfb2KP:&2=>S&6BV[-K>H=.?XQ6?<2
UAFedWY9aYI?>M]H-\/L&Z#-B+D#d:Vc-#8S.;31>])8+1^[H(1KU=43Q&f6ENN;
]#6(RR9TV@P6DRV.AVaY99W:RU.-=T8-.)-d<U15B=++(/<J&?7&/5QV22GH\Y^H
OT)9B?=c_QFU;)<b8eAeQJ0S;P;>97@D^?4=2c=1Q/+OJR::6GcJW@^d_aQSUH^8
(B557@^8G>H,L[&L&1B7PH997J&3gN&@B^=U\H:_0<g:R^IK:HOSR=OR_E5-6<+?
E(?B4_]]<L<Ib,<UP6IQCCAc9VJLD:M-GZLT0@I\NR9V4^C).VNG57_K:M&6dQFY
c.+9PX@bJ_@XV@U7/66IQI<);&dCG?1]<?f]:<f_@R>bN&_b<JNdK(_NWW0&Da+I
2A8?]_V9=QC&+[b?#E0.R#764PZ<c]M#a^M804ZFUe22<F&_-TH4&,L>FMN?+Qd&
&Qg\K:?-5+-N&1G9VDZ[Xda(R9NG5-e+[FH4b[(5PCb[LLR/d60YWIU]/GDHdd:H
S5dZEP4.9eJU##6:7F,1dMMN67Ca#;JgPaQ^.DVNI<,.Q4;2#\P<FeTP0K:-6#\=
@8LeT7SXY1:]QHR&d#@CLNQA#<-fY?5BEJ;[db;_DBV-H]c:<S_O7#YAQ,)^XEMP
;cM<>2\J2^H^-K<)6YdfS2O411ZHGSP4?Z\F9])(KR(#+N@IB5@DZagG_ML=MY-c
;B?+Bb-[_GJ#?I7C2X2^@JfT/EM^JP2CGXJ[JOA(QJ?#VV-+S85#KWGQ[36VGY&e
9[358;7S#W?0+)W<dd@:FZ/2(g+:PQ0.D7cY)Bb0XaA@QUA7J9(C)@;]AZM/ZX^I
L)O5aO#/.VR+H1)LZW@9G-ceI;L9a)JWV_8MD^/Y24:)PJI<5RVL@L:/#K+DU7Z0
6?b5_=8NK-:OX/<0/\K2;YY6QedBO3DRH]\]Xg97?7)eY?ICY5-QS4FT2>=0/Z,7
JOPIY0>bd7\g_#VD&&YH-eYAL/3I4/I>9KNBNT<[f#:Me>JQ90EcYf&LcN5=&WfI
R&U6CG3M-cRPQ)QA-6AMZ@(^cQ@(<Sf&5MY?:g#Z.N]:JR^X]:9R6++J^a31e[?B
XXa6MZM]NQEQ1AQL)NHYeXe\.H2_cD9bPd^@,\>1QbPA1KCAC&4<^#T@JJVJ;I&]
[<Lf1bAOaGMe:EV,c2_fc4D1ZHQFXSZ(/&]fD-9(SX(@C)N(>@d1&Z4NGT3]CX5f
.HZ#?=?T@N2O/&GKQH6gNNd^d4XeF.3W@P3fg\bgC]1+<_b+O,B1B#dAed<,0]-M
g[@;ZK5IQbK3PBI6QaV<7(4cO_G:<[2.1QWV.?S6Ge^DO[A]:+3\W7323dSL:?[J
6N>@C:^A3#H.QUWTaA8bC.84/.2Nd7SUCO^,6X5&SbQa;1TI;<QYbf-H@O?17?Y-
d3<-1K-^Y:[MDB,OJ:N]:U/TH5=c,:OM<_B6d1aR]4FFEW^TM[6aKQC/8L^D6OB0
gSBFJ)18(P=EVGJU?27.\8c+V,\9e\bgARbU&GPYSYgQD,4#KRZP;5ONc61;E+^N
A9GIU1EV+CJ>\J_=QC#7:;?,KMdSL:EB0MgLFWKPgX0T4UeCO&7AE0_?,PSZ+]WG
567UFL^7MPa_;A,>WU+/E^N4VAe(a:A:1^=J1eV>>TS8.-#d(Y,3ZFZ>1?aIS/+E
RW[_-U@P2P:f9A2&);8#;E(3g<4D^b>W^[Y;/\Sa0GY:L&1JX)e=fN4&_Yea5e6#
1[NG7UE4BD&[cfA&e;&Xe/1OX\)e7ZSBW_?L>QCH80/BEYNf_<IeM+8B/N<&N/@I
(^W[0-Z>NH5VacJ,#_CXJ>D-J[G7@.,UA_&Y+>.Yc>&/dR)3cMZO:#F8M\03CQ;R
8T/^DC=,6XTK7LOL8O&R./,g<Wc>Y@._G\P5V.=\J+K=JW?V5_4Z8U>LE3c;^Y-g
10#?<KQd6FL</VHL4QT?C-]R-?[gAgQ67V,S3bO.8Pbd?CE,5GfU/>:?0KDIVD^Q
QaJU,-[TLWXb[5MgU))c5[.30(645C(-P?eUM;CHTE<;D.be-<MgC94_FP)\]#<>
fgHNKZO^;4GR:L4bV]BTX<1Se)@B:.WJV7(4U2?M.XP-beSAMK/BB5G-g@IU,Y;g
2>Peg;P[U?7\5OB3L)fW@U/-EJI#3^bD4/Y?a9,aQ^UG0GWFX1X&K+UdWBABE<3J
1YNS^@-?U:2Hd3ER+UT+W4I^J0RPC=+eB7LK\9]0Y)CI(&PT]NXD(<cHIG12A0eY
C\P)V_5;P6,NRR;YV3=/SZPA634bT>-D]N^_YJ?:Fc#USN@)G[^AAT26Xg=IC+CC
F8?TW:6fI/cN2baa@AKaE+Ta1#=a5Z(Q,dX,CP/:6[eJ&aF9E0G9Ia,3<e9]g,VJ
-LdSe)8/Fg-QEg0fU5WH,TW<cCSU_&318OZ(:F40KFNU/9CM3f5U+]W-Y1:&\]T>
:V)?QBS+MG0;_dcPB\.QU4SWFT9PaI[c^,I(bQI>D/BD(Dc4Z.M:\7^N^4AQRJ1X
IDg@[5#5\/cJ3C<7eI3O\#0G^LF39,c_4JJ)FLfIN6UIT.#dP8^cP:f\GHRc&=dg
#\0Eg>C.\.0A.B?:1J3aBRE_/(cLa<F#+DN:E54C\>G.J^V6=[NEKSa\.eR3_EDM
&D4P(&dYU4&[fMWV(IN_\fK.+Y/51>9M2<JES)WPQCE[^)1\_:YG9F-LQYD[->C6
9?0]7(?K.D9N_H@W.]69Hc9dMg>]V3>>DL^IH>9CZcdI3HKLa0+BL@J_R1YMgN9c
Ac+b;U)]Ga/8WC=6Fe?8Yg^a#]PK\L\&?Y?V4_]aX+KDF(T>T@TO]M_^^J\.[+:&
Q/-@9PCgVa+HdJZc682&REBH[.9.9XH(JQV-(E?a,A3g+ILfMf1:F)4SaR<XX&a.
U?JC/LSY;.C/[S_f]ED3(T4F)P,[Zc;SVELD7beW\;E6_2c+2R0=)ROAWg=+AbV+
)+XIK8>43QJ6K32PbAIg:4P>\Y=-@0VL>1-DI2DMRPg?MdH582b9;:@KZb2CCF1C
B)&+eK+MLOcc,TM&KH>g\.HVVWf9(##MdI_81bS)7Q4DDS^K-55<^Yg2ZM&UB>K>
GDSaa=GCYT:&X1FC;:.b><CcVUS.S4_@0fcgO_\9X((QU?Q(e+:S/AE._HUf57-X
]/P@b3TTFVK07=UC<JbHMIEaNEB4:e61&gHKQ&[+\/9KbLT[U1NaXZH/8DPHA?d_
:CU@?5ROT??b7NbKGWD.YG(D#eTXN)LPW#=,(OTU&=NQEBPA4AY8c_^KFgS2R([G
a:MaPE>KY-8YNdOV39/1Dc4U?0A_Ac@:e.3&[aU,NI^IK^GZ4AKTNRM1VXD-SXNL
Mcd,I]dX#(5U)YfW/a_@/)B65LZG&V8D1?BJX@H9^PIa]T\;7ObUR\PGSX)=L89,
IDBB5F)RV)MLO<\IXScBG,<cbW?OZDCcQMR;[GA6_fQ5)(L0<U(=[@b^Wce-7.NX
00S=[6U3X8]UYXM(9<U8O/:@,_==(/WKeY?V&]_FFd-9&YIQdTDMII:DZI-4#_A4
>3U&GU=c8HcfU(?S8E)4,5[@SGc]:^&<ZQNUNFV==LI,dJ,6FeC&+F-])X9dC39U
69(?+9#E@gJZRKMTN<U_c<HRUaASaUA,(^G:=H9^9;,7O\&7B^XbdB+U\KCRV6P:
f9H@9+[0A-4;FK03dfRb\992e7/fM#2Tg,;>))MKC_c/@KXW)b6[Nb&J.#VReM=f
+ZQM]\A^1g?YKdB61Ib[29[NJ-:S:L+M)6W-(:@J)CDJcF6Z8R8/)9+87ZHKg/8+
&g&->E3d(&R4O-F]_K>T)_-[(&7?M4.&=1[/0<cX7[a5UZ&W0e=;)@9g07dM)F?U
.OBGX996R3#RH=K^HCM/BEaN3I^<6g_\W\1gdA,K:F&G)DW_-]/RIS4ENJG7QE]]
>I@M4E0TWD?GU8fb3VR^.F?@f<e6>X=Q5<KW0&TgDJ606/W,1cC:(JXF#9M<?DH/
CO;cb.?b<e8>&U[ce<R9.79H54YHRVOBJedK+UN60&<AQ6MP[.?gCJJ]K<f,P>7f
CROaWKK4VO9&YQ^VV4&g@9/554;7V=Bb4D8T0AHJY)PU.;U613-YPMf@e7f[44D5
gY83@98fG>.TA&A7e#^&Ug;g,E=eJ9Zd7&H:^CfJU]B>8+Kg5R;Zb#g]SKS#.S5L
X.4](]&M@Q0bD0dQRH;N.IU81\)__W-#(#G5d]DW9PVH2&YM]#cM]-L;RQ3LP0.B
,cQR5T-SCab,3IK2.DX/L9SBgFc^PAXQ\)FJA@]dc7,M9RVVJBV4g_?ae-VH#8(I
aXSF+T9LG<W0c75N^>\U<9>R47g)\:KNPKXU8):US6Q&PER<GZ03ZR><P7MeE&<_
:BMIe0O/5EVS7TV3)+e:6\fYL[GKW(8g+&B(/5^1KLX/,E]3H>E(:5cI6gGO@^9,
Q(GP<#Ga#X+;<YPb^9M(#H)^UeCNIZK=??A/)5)(YH&,CBAVIT+37<#W<QQP=6R3
:TJ(I11M,]?W3U]cJE#g)TW)cT3@;Ua]+H&Nf3.29FPB1)C=(./Y<(+G3^4XDGNW
=E[dCY[SJA5,aJdAfRB=gM0(_Y))A(<]eaTZU]LYeOE)6a(YIe>_MaC4GR4)eNa\
Z9GZ7+fRK^BK#?16>ac)QCAIO5f5QWgOB]]FUIc_E7GY0?V_EF)?\;=>S+4HX#@@
5&:ZgS2<^K&,PX3EX/g=FEXTN.P_#3]G7FW/X1.]dK&FA=A0QQB,CMOEE86<<8cE
DX9DH^;;<If^aBUf:Vb69F;f_F#6Y;D^)c<@KJ\cF<<^b@YV&UcaU?=.Ib0&1)ZT
Nd.6W3fK^I&R@,\I:_>GP:1KG1a/dVd4Z+)[[f7T7B&IP9Y&XW2g@;1aACW+^Y2a
&JNN^?c&&#T8\52/B9TD<M&EUIeO;Ua#JNg8]II9RRfH9],#f9Ze1ZE&L-6Y@>9b
:R,-dEH=8QSJSI6d.8&(IF]MPIU@2__W9B+&(ULRRd0<H#>G8JE&7g/dEg2eZH+^
9B[4;-GF\,JRC3)J)>5@_PE?fda0XAZZ,X:JU9BD.U&D^4:gBc=@9>Ec0FO,9AIc
&:O]&D,[>^MB6VQ[T)7eP46IVS4#OJ7ZIcYZaF;I+7WXFF[FML<Rg8ENOHU<\#:9
I7#[-^S-BR[\0&<,;-KbD?_\J;O3M,=L<1ZR4L#6Deb)CF^;_G2]aD>LFK#(F9[a
DC[g;C&=-E1)>SEBdYbb6f?-=RAPN<=GMK7R\L22/?(TC[J_@[1H<PM+D><4HfJa
>L/F&.6XbHT1A-6de:-U+];c&)JKI2Z\ATCY6fYM4Fb^d;8Y]@@ZT--f_,(Z8MZL
4J)HE@E\<(dK1L27QK\a^E<@EW4fW/):O1=00f/DfN8JMK2Y[-VBa8ZXX7AYeeS6
N4KSEA?K2/[>^fXN&Y?9f2/_OXBfGK8b,W.T/41:2LeRK(L59M5^W13,Ke[_PbZ\
HUSFST;:V@QWg2>1IB(Kd=\FVKbH2D75c(V)Q<](\=e)HJ]B7gW8#)Ld^YICOd^;
[MHG:f1Tgf7WUcMG[&G2Z&&]G).L12f)?B:AeaB2(W@^Uec?6HMdV4fcR&7a\1^+
_&f)IV^X]e)0CRa;.YPO:3X<g9\B26\(.gM?;#<08RPNMIa#+06MFTZA6G\>A_6N
2FZ=ROZ.dWE,Ve[^B5AeEA[AS?+S4,-)ME5P>K].+6L4@1),E>UF4K(3+/TY/1a3
V>(b:bW-375.VFC;gIM7NT)#</-0.<H]AB3fRYDSeJ&9@VQJ1]&O6=3e.(N<(EW+
+egE7-8N4Aeg;N;ZN:I,A-+NC4(D1?BM-=DVY.)aX@_Y3;THAQW.4fC_=f_1<&57
O^JS\_Id2VW4dZSUbM01bPRY[K4cXK\3CGY(b/MF^XS/fg:&[RW::.\#1MU+VA]Z
-W11#Q6]JLIdO\1]gU=FEJ2P;-g4=\@A4&^&-FJ]OKL@e,9#+.@aO=]0)782C4O)
#D@cFN,GN:A?dR_:#L@T8Ve53fVSNdX]KdFC):)@VX>ca82L35b4Q=R[[E51ZMUP
N_PE(IbVebfTa=eaQcbC?c3=E<,FM?AU,_&U5+/#WAH,a:eOP4JZ8+b3ITfH_U.<
N2-[U10^H;L8UYND@,EdZQG09SI&KMPaK]</C;SOR3V4R^c>Z>G5)WPW9&\,_V:>
HHe9BCB(W]@R;]@5B#@6B/LYT,5N7Te,d=M^FMV#7a(0\V/L(<I#9Fg?Q]F>_fA&
6;JTaBMc9CBX1+W.9HT8OF-@IQSN5^@)D#5O@]<4G-6C52NT2W?f+O@WJ4[9eNbQ
N64A/)C-K3E#BG,/2UA8d5B.WVH7S24];Ga^<I\@&5DYSAUJUe/NO?C^C\9QD>UG
<4Ia/12_PR_d--@KS:8-Uc.+Z9NN(,9CO.JI(:H,)^?/=ILDF-6a4A30CM[+MBHR
TXI:FJY#[.K3H\aW#gQN(TJfQ_.YQc:6>gEG-g].UHPK.#K=/[2>(I/,&UIO,b3X
7EV_7gYdA8Pd]Y+G8]ZeYWV=SQ7Q<(,Z\.Y7I3=7;=[@Pd;UWM\2I1=TPb(=@d>F
XM^d2c;4VWLC-PeDLZJf)4@;J#]L7eS/UK?&b];P,FLUT^<C=\PO6[EN^F7&HaIN
P)+<g\0cSEBRS#B?)88U@8QG\G?\D#RUL9.>+TIMO@ZBWe?67_U.-#0^eVM:\YK\
Z-_g>STaS+@)gO5gQ+:A5F&7bf#U[L9bQVNZK<ffLY[I7&g3dA2,T0;0@\X.\_N&
FEDPIT3/OZ=>fH4c/c1@:#,?GGRe1NAQJ&>8:.Ne#E.eX)=[@Gg7eF0]DJR82KbR
F<KBG&Q)P-TKYT5K@^FaN3#+CAE3Z?C4G4E.;IE11_LV;d:E8982fC+<3C^R8N(L
>P6b#@@#/c.]L?H?U>d5;WXH>.cWYO9TP,9SAPDCdG:=R\BSQOS:T(FCG()^T4ZX
X]@e#)G\R_47\9:.T\MI3;HD5@L8@7RL@W>/,^))FNP#cdcFd4^H\DP)2,cVHPdC
6XTYY1H>^K=<XRRLQVTGf&cMV,[RSaO@EL1B<YNB847NaeS+DD,>R#aA]FH/+a:M
CeEJ1c:B(IYQE]0K0VCOcEI8^@f@<[^@.DA5&A<a;,QHaPA(d:b6.9<E0@&BD&.a
I(B:=Z4>-5I&5.9337TP9fWgf,bc3JQDLTfN@8YCOg74XU:_JNCg@,JaN9L3ZcV6
[C7B7:MQ8U@g3eM>YNSC)YK-JP/;DE@]V]X6>I_9BMH5+6O/B2DOL^\V1B0C.PBH
A.>H1LWf(8,:E+a2Z3f3WEXa<)S33]?@(JQ0KOcc#1+-gOf4;(JPY?54\+(LDbFD
G:F,7?3-.eYP?3<c@;XU+e,.(TYWU6?X(6G/LBbL+LIC&-^G@/8WUU]5]9:VQ]#.
SPHZd2Je)4G+#\J#P[Xg40_\P)T#JUSf\3dAf^W&L-=+5YJfO0&[K4T@V\a(bIN+
YE0-PbKNeP\:b.UNJ4>81Y[-I;^X?#-F.bPW<X/@HdEYaA<#7LEEY8=7X5;fKa7=
5S[@<92NS&Q?#4d6:@e^:-.M7NFX8Z#5GT6g+NE(4CL/bF5#<eFfEG+WdWB5_VCQ
7F:A8>E59\USL(P4g/P]SP^^U(5LH_f+F0e_e#(GG?YZGK/<^VORNcEZH@#e1Waf
&gZW]-AW#2T-9AR5HYJ[;WaEYWESTe.M_]M\:2WIc16=GA:DGdWE0P03BW>,.UXe
2;?6\G/6LOfFN7@=;I0KSEX(RI1P-4_POb37WQ)F[>M;VeIRKc<73?ZFIIg(,1PN
[56XK55^^Q88aBF)JgM\\TgG[K:WdbI2/?b[KX=RdbHA/>]SK&D)_egX#B_70(.6
6W2_\bYI/2@OPA-^8;=;9V(E6+9@1NYe]UWQ+>/O^8B;J73R)B.f-R_F0[WLeLS.
E@c;4--NXG:<OWM4DLQ+_IE>,2Ca-JN19=ZJ&^#YOR4;JE6b]O8^K=c.gEZI_9d\
TXZdS<JL(+Rf4>[+b#ffe>?&;>^AA5bN2=A)LZ00SKG-[?JZ^LCM,1^TC>(FQ=dE
\2[<7K</#N>gENEQ_aH+FE.@ge@81N?eIPGE7@\0E\PBgEg,FUS?K_G4@KPZPQ,)
D1;FH,be^DG7K;8N=OXX=;e5<cH/[_B1T\R9)FP@+.A.Ga3-NL.?0+S_\>;SO&J-
P\R.=eP2QTd_(=,?d/9O==S-=+CB7BD.c?Q<0&#Q+9FD-0>=AHA:)NL--1S0=[=]
3?);eTV],8FRLP4-dXT3gT63<JaZ=2=B2F#DT\^._;:?=Ye.1Q:4SV.<SPeY)\I^
R6K(EQb^T7L;5P;9cAYD@;bbCB(1e<U0++GSBR1g=f(ME)3fI)1f@0^QV-AO./EL
^7D7\Z>UQM8Z^;JHAH1&2B_BG#F=UYC\Y6U[aGQ&O#4=>#FaWd>Q=#^-WW3CI3Wb
Vc0<^LI/gM@U:(MHc(@VG7#S\=4?+CM61bUW3ZK5g[JacS:;[5^AcC6gX;H[7=d@
O/OB?Y_g@)N6_,e[2dddT&\=f9/CR4U=_1:T8f30]P7IfL_^7>8Z16A9#]?N]&[f
U>X/:E-708BJJGE-30&S)7DeNX8MadTdQ15SUg)HXWD9#HG#S=cBC^3RCG@\>)1c
8aM&X1UMdeEAM:U][:<G_4TU]<B0@cf116DP8&FO_Bf9+c17a\e^edY<5eV:_71I
8<?DJA<A_<P5LSZc.fQ]^b;)Q5P]JX[/a^.cDN0Q()=8eG-S,DeEGCKUQT>b&d).
>eD<3;+?(b]DD:JP##0+(dNG9U-73R6A\X</KCX;S/LYa[aUF3DAHJE93VN;XWf[
VN-;O<<^93dT&CN]Ycge#S(0DKPg#cP,.N+M>O8_==[>]3@//FI9E(+WMWOJC8,Q
^cG<)54U2N-?4CaMab&#DK>BE1(_&C&+GNH,TOKc(3UdT;PFVSCCf?JNL6#9.VN+
,DR;YP9?N?@AP@VK#b;bVZ&_/Wb])W<AQ>UY,-N[:HP5+IE?+_:_>OJ6Y+YGb?bc
0J4)#]>4X@)L&EC/Ta<fL@;-ARbKU#TH8)A+aDfUa/6&g8X[MY_D6P6b>-@/BTQ1
c>E</4G\WZ0bZ>:a^g0^SCVE4H&8f\Q.7X1_+,^?MOY.Y24[?9[+c?a&TD<,3aHA
#U&E45RYg03ccg<(SY>DS;379;cX9d;UVBT5QMEI-GEQ/D(<9Nf=FN2==,Yf(U\5
3DQI\7GeYZIK.1Q:f^)5DgUI[P7WTSG^dT2F@W[419A?T?R&(](<J(>8(+QN5F=^
&P@X;V0:P>Kd>TVgV+@4Nb,=APNcNb1J-7ZS_&(2^cNN7?gJAa.ScHL1SMOEX\R[
DJ5a>b;OX]0a5ER/L^5cgVN6g-4F/I3G2J+._F=#GaOL?XeTBH?5@dI4cI+^;A7g
Hc5U3G>5PU62<[:]5V=>WMAP[0W(M6<Zg5e\)(4V)M&EP1L0?cSN9XXLd/8(WdR2
J;23,\&0[ZZ0UXdUFT)9M)EC=:e+_2R]c5[Z9+;DKH9IRSA7+<_@=]]OXf:a1D&E
La.eC#E2Mb7@a\?;:R9[5f1?+eX9\-QEaUN.\QI-NYR7EPZe8UI):N,WFbZFa7dK
)LW<73-6MM&TAAXeVgeAMAAX[[W#K)E1e@gGO?Oa72\f-]f&HAbPP8U#[Rbag4^X
@a22DVWUWLOLX^DO26+b(,#cK[W_cO+(<5;G0G30UQV4N?:+\@TG&TTHYH<34^F)
+->JX-4F@?/7FVGH:+GR3#e#I&I0_I&NbSP,]S]8dc7WBd.3_]PGcH25-Y,]07VV
/WX>4VX4BI?dNG_2KA3P,[YS4:BX7?M328[RE<HK[H\2V6Ve:O/SX_3dTJFCOR\+
M]9e>?9DO3gA(/VG&8NLY.+FEQgL>+F6>[4O2_6GR?H.U8T8HEHcA1(cB_,UZcZ6
MP>#3HJH;FZ.NV8:b?XYLeXTC-91\2N?=#NYR,R)>YMP1P3@:Tbg02Y/bJ+-[9NO
Y=_HC=f(6g]NKU@?]QQU<ESCD/#X+1BWB8&X@7.^>ZdW-3_gD_IFBO0G^\##043/
:,3U+aKY;8[0&7:0LX:?MZWT<=V7I4Q=D1YM1HV60X>].Z?99QXP6/?\gX2.g@fa
CO7?aYQA<,EN(d&@6Y)=+=c9<9I0d.NB;M39S-I:T+=EA6CCK4L.gXA<C3./dPSO
R1a5U(_(X33++af&QZW7U;9fXD#HI,I8d+[6:[?S+#,7WS2Q8GVI,+(7R:I@0#<b
dEOQg@/AeBNN_J8g>B?gPV[c)OZHBR:R9c,BR&]G;MKZM_SHVX=L32ZI\USBgSS+
(BV8BeF1UZOgKB)(MRRZ0EZGe-?L0UR[2S+?<\GKO>_=-T:<3D]8f7;b+f&5Y@Sb
M/dcK7[XBC1-/#93gV_f0S0VLR(4?dAXB-5OJFMa_1H]\F<J-)X2]Y>#Ub-Jc?,V
0PA4C;0PCI+DH,L64c[#_W0B6ae;5P(HSb)YZB1M&59-3(&g1R9fEe3;ST:T&1AH
e2=/REQ<cD^]OT+Dab\?Ig@]=5b)cWJXQ9P1G4Z5FLc;W--8S\9)[R@II1\M=bQO
:UE;RF40;[BUW3C\I0gfZ>cFHB=]B>&,;40KHHf,-PA6@;K?47[O^2,3QM506:6c
F&Y/dG@fae(2A@M[_YXS_L+=c]cGa;L?JU>M6OBXVM(c8H4C:7L8[CSZR12+Dc2T
)/],-D0?eH]CWf4[ZFYY9T?_\89TNJ0B)SRJ&(.]U^UFXLG(&5<TW<F3LA<dgPN)
/K)#509QdfXCY,NeIdKg1+gZ09IdPMf@-YWT=\ZKYT))G,.EE:OQ\0A8T^.\K\_5
#EC+O\.ZJ[B=7PRA3BWLS4<91NN7)(G37:/aKH8D)L,;P]=/0Ae3T3a292e\<;V=
4+:&A4XL#SWWCZ1G48DX(3;];^L2fFKOTc]=TI?L(L/#N.OEK=Hd8TMe[_Q1]fVD
]2M.Ab[[ICDeSEc?,CNU?aeW<G2_RdR9-4AB8Y^6?B;W44eS28Ye\2G[DJ[NRbT<
>7[-)a<<=#A/a>NDabIA?f4&RVC;6GMB<GBY)92H\g,0/7J[#RBNH^-?)D7V<[B(
P/AX3@g<)ETTa.HB6(>^3g67MVRCOR=+d_MDd0d..&QPSZJ;I^//^8CH6()VUeTf
fc>>Y9\-+7dT5FC:d7PW0H-15#<YgO)M4bd@4dHOZO8<1+;XQI-2f_>eeOI+S<J?
.L+9\IIaaX[BQD.<9:Y]=H/R\;=2Af?.X>g,\d]a30GcY59PBfWTTRZX>8LW#8FP
b9Z9M1,f=3EU#9c,eSVU78LY\XJ_3Q,G>GfUV]0U\b13?Q,BY/96H\.&+R/69/JG
\ZX&J@bXG((?PJQUH5Xe^TXMO05XFR_N\<_X\XA-8WD2:ZG7]W9E(,;I2A,IBdaL
+N>RW7F&HEPU&(/da@Y&4@?7W;E6De>8<#J<UcMB.b-aWAIIGJE9]H,,d7dW3;f]
ea+WIf/BRUJf()-9NdGUZ2:XUHZOa)0=_Yb8C[OXDfSXd)^ce:GVd2H2E6cOB\R5
SUBFf?-M/B862GBc8H5DL<+?Og5)3CT.dPA1gb/8UA]JZ5AfgLKP?R[CFgU4^/[&
7J><,)RG>e3TJ:F13H5):50J]>E-^9Eg[7@c\fK)5TZcGdY0:>\7^cL&H<M_1O.^
3?U[P.X#;)Zf/[gDGIMg^J]eJ0).IZUd,,<M?H#5(_X+CX)@0R#c)1VJLb+\F,,<
54V6bMW=BKNARea^R<D&@EA,Y>VOZ?WJeDE@]c\^9^:eD=N1JAgfb7-.+Q.B?/^Y
U6=H\V]R::>A+=L#<QZ@5QX52QS_D&\@-BRS9c&Ab/4Q:>0[fY]#.D+3>?#]9KXL
1-;SIC\AgQE^,MBFOK=.J,^I.f5:.T_2YTG@.\aDF=c@76K#,0?&&UM4;F^^JI4D
WW#]=#B,@?<Y^,PEG8(54G5OgYY\6)[..:OEe+UbcIC;V8RY:Sd82GEF2>[\\1N^
3ga.a4Q3]1PEVWgR[fE/@USLYIX=JZ45J(@#\[D-N&J,5&;9Te62/^7&(/Hf.;78
We.fT@E](4[KB^S+?CQI;gb1S&5F]/>@TJ,:PNLTe9CbDWKNZ;+cDXFR8AWDN/8#
Ld[R,P6G=2BMU^^7.SKQK&(=1c\d[N>-H3OAB>Ac[Y<F,Y31I@>@;,51O__P_BX+
2KQ:\\fI0C;FP(347X<gF;+]Z7DbfT<f>D;6b.A?aPUQ(X];.M<2[&H9D#ggM^M8
4bbG))f>b/\B^d0A1,.)Y@B<IZAZY0\XMV;a,V7).Vfga(e)(e<+ZCK<DYa;Zff0
KJf;gO4<B<+DLfbX;U/N.TK_<G_RbML8NNL11NSR@2=cW>1L5&f-O92D]YFaOWM&
/6?^LAR<DZ3MDKg3(BG)&M=bS0^O:gIC63.e[,BK=f&<J1W_;90QBD]5aQ#KN,>;
/EgH7c_R[0<[e+^Bc64#W1cKKX)BM^B;7\WGDNY1cT:+2U<MF9Add-\c;[f46d8/
dd4#C\3^F5W:C^DI?P[Xf7<32<>^Fg8D:TQ(53CB-&MP,);.9^DRY):0S/_1CZHH
b1.3TEa/-4P>+_>;dDFeF/EFCS_HE2?BQ/2T?H([d8WL/O@[KQ>FVg1621I56L8b
LY[7Xd7a>4H1\M/QD<D;(<&0,fO)0@3bG:dXHKCd-^a0J3OJ@1=+&IO-<5@U.CWV
7?:5T>abPZgb>;aPEZP@-dUTRRKRJ(\_8YfZ]?;7>KK-]WGV]=&D^?FgE;.7E.N0
UY(\@_^^6b85b1+Zb:O@V_M/_SQQ5NWK/\LOE?U=L/<Vg(Z/I>XG^87\?7FWUU?b
a>-a1J8CWDa8GAcN#5]A3W;IO5JX_O<[dNHK&:R0V4/;:abRU-GLEU;VP>bQK,K(
9.7C\<XSf_+#^3Hc1dTUAeT5Td@e;G5#TX^8?25NR:Yd1?.8J8F8HE,#(VDg,<NW
dP7(PfULg6)>J]S(2ZS+H9WUdN7Cg?ePAfT(K#AP@X#WJ/fP_Z8:+D7YYL.g)/1V
\8\4?2+,ZJTUXYI@Q=<_Ob=7F035W=:&6Tf4=<O0.IT;6<:&L)IVDIZD+8JDE=I[
f0&U)S/SCE>0_IeK>#?5JT5.(KT3Q-]14aR4,5<(3U(<K.0(@aV:00#:^TTa5PVD
;=eJG6Z03FF57O=GN.57VM4B6:QJHd(=K9_f5J)IWe_eA8aE9dQ0GE+G(C,dFOYY
4fG,@cH3H4WN:YgT0;gD3M@O[aYeH[2LD_8&YY822U,[/SW7L#Bc\G1TBcQP7@IQ
X^K1/<a_5GQ9BIB8EcNKVKDbC7?)gLG:bJT9PF333DJYUQ6,Z/QIe2OS/<SO^I__
4.<e2.25][K7S4.GKcf4b=:10.&,+I3LW)RJT<^4SE^a5cV[8(.;0D;BU16=[M4&
AUE5f_+-DdJ=[TBFcCa[YEP3MgQD=;/19=MZ279PKE2VGKa\[Pa_748b<Pf,VC3J
[6_V>\UHALPP9e3)=WPL5LWecD:ZCI>@AOad1G8=Q3WL;X(fT5)0IMaVcM:fDRJa
eYF/SP1Zb?2I@W89,53Cc(#7VS<U99,#[+;UT_^R03PBG4<7d)bRgb<F\=DgfE;Q
1Ee-X[B4XX2.9MGAS<VCR^)3c(\eCVCeIK:U7Z:_afX>bf9/BP0A,LU_W6)FK>5;
QL318N?+K(da-.DMQcXRZQ#7@.dW4DJX_XI]-]Q3ZONa:L#gc+MVL\d]JbSTMTVR
&-)e71E?Za6-1:Y/cV1HP:Rb#<05A[P(#8A5?Y.N]P1S/.3=1d3Rc(0-,ZT-d[O?
b3]5/+D4W9d<.\fN;VMX_WI;2/<7&[WPY3L>Y2GZ\.eDL0>W\P0Ne?;?ef&.4&>8
M9_=<P9#08Q#X9VFRd_OF_<fecCfMEa_3KK21Z^aX\V([-_(3NSSALE&NMPU,S[E
CJ+HI6e_.HE57_CB3=>b;GPa9aSZ6;B;M+N<=^._,(3KgX^.SJF(f:YQ\#36SEZU
<NU2ReAg^ILC7IO_e-L]0Fa(W[P-dX4#;0U2@b\LP;-A,&#,-VC0L/Zgd\>E7G6T
RCSAVG19Z:d__49.8eKEd;-d^WbZ:+WXMG<,ggL,HTN_-#0d:K4_a46b;=(Z12UR
YUWVA>bSMgcKI_]IY:)AaL2#[(YJG)5>89M240Y>8g^ZHW1GC2R\#dRZ2DWMBV+&
J44YBNag?0bHVfQV2>CUEKC8a+@#c+e>719(9,\Le+6L;6U2@6dX/8&0H?Jec_bB
g(9U#5dXL1T50^UE4cf)YeQ)L9SQVU?+BWPO9(?2,7W(K-cPgf3AUaSS4Jf]Q6J5
bSWg0_#P39YTcG.X(SMAN?gdN1<MXg3Sf&;V70V:e+A:ddSbT-\WN9L>.,U^;3M5
FE[Jc-;[QELLf460[Z<?0W.GM(RgbfT]d&;9/G32]aNQKR@FX;-g5PFF.>Id=J_,
47ee>(fb<.Ce<C0TZ@cJ[:Eg+/X:8E#c[EZ]1-.=G(]Q#LNC,</1S\]G7[+.aSBg
O-(44P9ObBd\ZWA9eJ>VV@)U2>_7JWMKN_)9U>.\6=8K]KU[C57J@,AD97e=d9XD
,[VJ(NDX9>=6(K4VR)G\/eaWH-TI8ZJIIRUbI2R#.M14c3]cbJ[3NG+L^A8d)QQ.
7+RN([?FM+AAH<^#JY^9L0H@AHf<ef8O3-8W9^HX.K3AL]314I6eD/,@Q@9VJ5^Q
(TKER,abOg&-I4a38;MC)MX>;Le;<X#a6c2Q=^RYN^G>/I.4LIaU[d9?4BbL@JSf
)eBfX6dSb\&Gf?,;-WUI3:-3gKOX1)]DQ3gacA&db^-C3g>+_>17WP3c)ON@2g2:
T.05<8#[W62.P&7SM^^_=B4O9YE.MgK^#ENdF3U+/[,_C#&/&[S;A\K/@/BY/D^b
_gf[&)D:Q11<J\,B?X<aB,@NJ)EOMA50L9V>J#Aa3T&WfX.QSW/dR\)e-)61R0(2
aG2T(V&;J<OF7E6bXH@OKI5K_J<+?VIeFQIQHQ4TKHgAY&I;\[e>_&#BDNN[OMU>
8?#<^^B3RKE-4_#B)3BX:d5dSA,=[bW<-0Q5>>ebc@L;d3f1<\O/dI#]e&d?c.D8
BF3H&Z:F+KQ@)=#9YY+H\QYILfg)A=X;I^JK#3a&&[\SFS8(eH#eC.&OSRQD=5OR
0,C3?43+]FX<XGfY84Z5U?-9.S#T3EA&FaK\cQ.a^D\@7PbL(7Od07=GN4::RJ0D
=a3I4Ye->ZL5OLVMaK9Ub_(1b[5V@FBW#a#\&cCE]cR;R69g/W3HJW<LY@QJf+FM
(\9^MQZ_2\\LKS,aKAFe5e1-)/dB8EQ<972A-2:Z#)d8>T40eU9O\[;LN\0g>b.c
+\,EB>N1F>L1fV)HI^g7CbR:]6dTC]e7-/)P^GEe+Q]L5=.)Ya\71ag7M.[J#5AD
#F?3==+R7IDH)Z\TBN]b4]0-D/^E^GARfdPZSE#A;#::#^A9;>74,ce4CD<FF0UF
)A/[PHc]2U7UX=BEJ[ZI11;18OP0R@FAK?f:XgdGG&S4ALfBVM^aB^UY+M^1(LWK
9A44N0>[3<,BSPT/TI8HdS1MOM3+JA793]R;G)b1SHbA#WgMY^,_9-Q?/EY<T:+0
HDS\;_Vc@dGY/)+RO1^8Q;.F4g/^K5&abB+K,D)^H8Mc]gI+TE[B,BY(GA1GdP]6
=@8(CGg2d]5?Z@ZJ;@[#:3@(d?]B)^-W0TYW9(2M4R^E;IM7bZ1K+EB@dYK]bM/T
>R:F7F(PF)I,)g8>.XP3deIS7[3:)U64Tg9#Z90BS4JI,Pf,:4e3-;&+GC3K-P,]
F_TZaNbLQ/gf?cQ6T(/Z=:N@0:)3SOY4@PbMH8CIZ3EebbCVJd;e#X_5PY;.\PSL
O?[^;JS(>Ha:LD5,)&cFUU;<=UWSEL1+J-.XW^ECZ#aS5@,4&<[Aac3;&P](^<Q2
75Tf=FbNLcUD0/PTD#M86ZR.VH\@A)LQ-Qaa#H+f4+^4bIcSC#>U.B43@DDaX-U,
3L?40c9#7L(:YSeee;_BTHPBXNQI,E<+(1P#V\W&Q6PHRCM\(\FQ]GVe?b#_GMDF
25F.8RKe>Cf/<=JaGX8cX2BgTfS6Gb.T#_=bVDO6K7GC#?E\/e/?B[??II2+_]8<
:OI-L1JB1D84[3EQ2N:MaV>(JA0:VJ;V69Q.E#33>#5ObFYQ5DL-C9SZ8YKf;OUW
(c=#Y3G\EYF[-BXaeGc0d&3]=F#>G:4+OWK<<Q(fQ&\M)a>Q^EOg1<GE(1B,8S6Z
K60:AJg=@)V7e>cH5NQ-=>cb&=eAA7<c6&F#0d:68?C)Z(Z<2=/b?3=1dJU.[LSB
L^:aP>J5JNPB@VTM.dB=@E,0gPBFYSRg].gdM6a-cc1WDH\#+e=a@fCS\-AdT9Fc
CU:KV/X:C1)PId);HX5B3RY_VQH4H+[7V)@G=?(B<7K-@4(>&1b&??8Tf9K>/)NS
#:]D(SP#4AV^1<^S(aK\0K28.f37GKT1Y-;GQ_#].8,H81d]U:_9e=8OU2eP(R@R
Fa50>0+ZE>\)G(VQ3+P\XQGRI+QaXYb3ZD1[H8XM#/_CRA^N[PRa0f^E1a9^HH:E
>OMI=TR3IQ(^5)bc.=66T4@9=C&UMb>9+[NDR@(TY+\cCZf6.P=Z6=K<Z6\eJ0BM
E[RZE)(;SQJF<aUD+5B-]ET^GWaMcgC&]V-8<e,^Xc[S3B8SE-HgGBb]9aI7.PeK
\D.BeLX@SYZ?dfTb@I_Ref85dC9]W3LXT9OdFHY+(28=D.3E2=QM,4cQ#7-T]0<I
[/0C==[>GHQSb]40H6T<]&>I/XJ#7^(cKW&<IJ>;@QK@.RfEU<G]Acd=VdG(K\Y&
-A(L,cePJQ-\_#V31;@O_A[_^g(Tf?#H8O)]J4;><Z3Kd20VL>Q\ZcKNE3c45ePX
H3^U7=<U3Z>d56R+J_U_FF0I:4((R\XL0(N4YZ,fDZce\,+NXRZ\M_:@BQ&/a.(3
-9@caP_U1/YM0[M2Peac-\gI>6MG=;I)_3M-e&B>GY9I80PadQDg3[8@:&503C/c
-a2G#N7dZZ[2Z@LEJS)N?U:2Qc:R;f-bOP/d=3PHMAI-eL/aK36dBb-0He\,YM?H
S@&:6C)f3bSEM;;1e6EX&e;)Hg6a<)Hg.ZH]0/PN]LU>bLHX0O,b]0W2&B@J1O+A
H8[a&I^V3KPQ9WFWcD#dQD/C_N6Ce-PN\eJKL?.QY)QT8F2@27^A+<4SKTeSXHIO
<C^FG:;cCIRK7:F^\#0:DVUOGW26UcQe+PLPR3F5BE,3<g2FgKfS6\.-#Hc\O-Qd
H8Q,WNXXR=G+3+6>S_]BMO?RB-Oe-+<#4T;LW[g6MKGESF[::2C\Z.RP?C@Ce0[W
87C,F1]b?=Qc1gUKY1;b7NP7@WCFf0-R6]4Y\c-Z&K#Q8DCTO\>Fb,9U<d#C^>(g
]=36\(;g[<a\R#]>7FA;^?^T+c38]2F=/S)1FE0PL_,FfA96F?DZ^<:KA#D6CTK)
IMg:Z<Z[P^OP22)T^==H:YGXMfc9@1)3X1O9<EDXI6Ec@(NfW[#OWV2UgW\)715&
c>^1XIDD?6=_WS_-#<LaU2CB6W8+A\VUc]\[WZaU,9aBaeG7L#^U@,(7UF[gG(;C
K2@,2_]D\))P?<g,6X6MI@)FW>aQa=7cCXU<R=1e/I]g0HX[M,f1?YBM3dc;PFMD
&QgST+PFdBf9b?N\U8G^G/a0e/9[64fd/dQ:fW^4L<\(-X)9^Z[AC]4#a>dWbR_S
g^)K3JN7F\F;\C:3#[f-:b-B)=G=/HT5D944]N+>W>&0E/XU\Y0IU=BCZ:fU4WdS
:(6M?@gT,DU5&.#LGA\IJ7](:Y2\IUFV?_4IYGVg0_3Zg-&4eS^],eS);0CQBB]B
V7&_?XdcLZ1RQEfR[;CM&+XLB?fE_U8N:47]9KX?:,LbRS9eZ5^O7H5HbSAX3JAc
=ANMSY@7@ELdH:U1/gL4N6]UH];<dTWY.VFO89]<BA,@&Q8+UAN9(&GgBIO_FDe?
F<A<QFENe+I2&G)9E#HQE;PBOI_]P4G5AcKR/_2T^AR?QNXY;_O3eR:3XcGf&Yge
LQJd(V\fKW@,JZ0YFNc#@AGMD_L5#I+cd5L/9_;-,1;Q+S-g7D:094ZCRJ5D.f-;
>d0Z0]IFL@I+ED6C>60Xf=HMfTIgPW^@#3d/9D81eD.)fb5^NPCI5OK4-#XU@ZQ1
O?Q;/^)8U3D6O@,5S(\MabM(VQZGUa;>.EU4P<cSUW\EHE0,X18L18\@gN.@<@0H
X8P\UXgM?_b8[N3)b):[8E.^2&&D2C]>Y+c-=8L5FC7A0^,Y[Qd]Q\>W3S)6-:37
CD^e.I(,A5&,+GGc)YH])V<f/c?(8^QJ;JQ7)?N]>f]YaeO:\O4(26=)3J:LFO#<
g2LU?/O(OD,R:C\+YeY13)DP+2DS,BZ^SD\W/I9=:-C7d//f6HR)+gQ.PQ[YD#.7
B]===L\NX_gBFaXCD,E)-GIa2cQOZ@d\UZ/I445(J+d[SCI9[#8ET@B]2C+;9,f&
,2cW=A/^:2=2d)R)IP.X,[4b05]Jg;3ZZeea1P@#KZQ-PF^T1f63#a=KK=bO+]5\
00DT[>6W-[F0;Y]7CV:.9E1UFYOL]H:MZ1S[M<)aC^9fI/2^N8B.e/BA_fP)]J0P
PCb]S2O/f>H.VP28acHGY3d<7N@M-]+N6708M(MCd]M8D2@UWK<=#&cR+>fADI.?
C]EYJ8;XeNAM1N=ER1X&1USVGH:Y&7a(>Oc=2MIM8\aB3#M0aNI&.,+]7UP]YJ2J
Q46[+#2@/TI_(VM3<DdHc860^,45\M8Te.E<<5)6GU7L+/6@N6)Z+-aaYda7[C&@
;U5C3a=e4SQ9K^OOH8ed=T-5+303[VT7KD#RE>]9)gR0[/7^FAc-GC#Cg3g4F5/:
A((;:Z64)QRR5F&\WN@?#I]9;afMKI]6F4/>2Lf0ccJ@Nfg2[LJKfQ#7E)-/AaA@
C]9XF>;2c]LH:-0MXUe+)XaBb;3/&XVfPd[5(]2/UHcJ331QfW>?@TeA#JIBC9[Y
_N@V.eYPME1H65/@1\P3TXYOWPfQD2\cM@D/-(B\6\G0]V4(_D8L]1#bD/gJMW_N
E_0@FE=CaU[Z9ZIWd#;VXHLU=R//85bbF3US5SNc_.IIB7G>bP>Y:^NV0;EXVO<X
G]JL/-V;N)6+Y#CZ^-.B+UK))GNNGKNAfU&Q)YQY(,HD0QV#bd65Q.0=RPfT0a6b
(1L@]@G[WQ#a)4\+RYD6[Y6NS0&G1HX5US.[F3TH2=6OT5,?&(dSR<QOdgCA4gI#
I,DaTORf7\(R,B^BA+]bKNP36.?\5]]_@M/1KLZ(GYI0Cf9H;&#&L;62eU@]TY5:
2O:/(2SU/IDD;5S>HQ3G_6:Uc/#_DR,EAYd/Rc5c8-U&FcI4_?8c?A>Jc5gC3Q]<
-:99>XXMF?KA2A;aUF2@ZA9g7Q<+E(g3cQ.gYRRQK6WFad+21C9\^V_7>+6D2XH&
3>>E;QdF3T\M+&Z=8=VJH(Yb=H^7^9G[]TS54M=[GYSZfV]>CN3@e:2PAe)(a/@;
9AF-C\6XaZ,7<:C>g75;+ZGJWARfOJeZI](.<1(G-I57S67C/8-I=J+29FMZdOYQ
B+DT]Sg+<<;K]V27?DFMeP;5bX0e/:073gKeI.U)54R+>cLaE;c7Ob+A^TGJgPLI
a/XI@Dg3J7&JE2b_Z9MXbgGI[97UN:8dH#^X;1D[+;P7@(V#&PWTW#gR=>g:bEeI
A[M@9f-cDS]c3LS5G?B4+-2)<:#Ld9[^M1+eEfXZT-3.&gg1]2C/&9B^A?UcHH)d
KR32;N9@NL=HZ3;eW()<AeO#,<[a7:<c9JgR3<<L(W]RB,.Q(#M[6Z5^HCGfTEcF
V[91S8@10C_I<BL\]9GJg1B9,4QP]T,AQDF_[8LXc#.07Y^cKAX>cPP2O,g(bU?#
^Y1\3?X5OQD:3bS/KACM2a8dd&0[-0\:UR2PVUU+0f>L9F7ASPL\=c3e[J4YeRNP
fK>Sc\[Fea8^&Z7]C3=Je6P)?.a26EBHMV?J,CX2+4<?49Wd=K[K<QO=KHVW69W_
Vd[G(EY(Z@_^V0?>&DMge()<1B3[cXGBZB?9T=QI^<_a(.,_@58-K(Q@)>XLPg28
cQ]Q6c.C\)61eF>F&#3cDW,<O-E5XB66?\F6;QW<4EF(^UNIS(cOHY=EWF:\1Y_c
P:,Y6RYS2-<#2-O1)L1c8LU\\0O.4NHT,<gB)AV[5)^b,6g_)e:<@&ZG2^K,F^6Y
;;B7+HYO-.+LK/+1)6;RR3,c-)#c+Hc/NO\OB2V9&F+4E@MaG2/P_UW(<\+[9]]M
dD<a3TLO?\LEREgg1^P0?1A?B5ROX(7:5&/)F_HBF1,f\HKS#S]X&M+HE:eF8FH.
^/W<?fZN;7G5dgL;>[cW2<+?W=&VdfXT)f6FL^a([8FCKTTRN[dB\5gN,IZ5DPa\
TWP+)&2^WS<UZ^IIB4=.DBU.YX2^.R:M>(cU>b80eZ8LOMN/=\&=#F-b5f;G19>]
;3H=6##UO4XMU\XbD2DVQ\-2AHQ#YI.>?>)<+Rc9cJ.H#f([;;,&\Q6#.V@YEGUH
aZUAV5&I9XZD&Sb70>.-XV814BW;@#FF8ZcPO@Z:OAK+CRF_I]=;MJ&.H_O#Pb8-
fPG@WF/BWB77SL:=e(^S<RX7d]B;NU;T8AB6I-AK<I?3.6.TLUY7G7f#Lcbf5GHW
;=59UTH?:TGNFgMM:fMXWJW\MOfAA3QG1U//[MVMI+@XTF7f-gH=Z&?DD@_cW)QN
TP<E39Gd&;^b60Le,AO@MCT+c5gO9N-,V:+0Ifcb/^[/eP5WZdIWD]N[eA?VM#(,
/1C2UeR&5ZU&KT0@C^579L.dWI:YOG.\O1MSbX2Ba12UCLL)JPY/R>Yb>V6BMGJ8
)d4)_.OI_P?KS#0cKBK:2Ea5;/eJQLV_J.=M-DcX@c&2@NVFf#g-4O;_6--=W5A8
b1V@&@/B0D?_WI,^_(2M29EEXNUVN.93GS^NA:]aSe7YEe3:\b/4)F-5WX&EM+;=
^S1a2H;ZP0/4:QLNB[@A+W5QPdO//.#4=Y77f+aB2OZ@+(U;MNd8F]_/>LR)RQ<7
UH6,X<.LWeg&]X,FR518>7+SK#5#[\UU3^MWQA8E&N\<d(F&-\EbV51K8I0OgV=T
4d.b1DPDVW<<JRT3AGS;e3P_1ACKEB\^EA5c/QK@:J>E4dXM^P@I>KHeR9D-(/@5
:(+-CW2Y0.9Y<_\EJPFO_76<5RM7WH)A)^:;5\A2g,:5EW6ZAg+eJ@+D<&2@cYZW
>-.>fcO>JKFcf_@3Z?>[9>?,Y;NPS3TJfF9:P+YY:IL<XP+^WHc/P2S@0+L7=&[Z
:,SPLL<HfAfL[=EPZSdVfP-A(7JJ(6T7f=R+QQ21L0#;;>5X\cJ0)9TRgA>bT5e8
Kf@Ad;O_Pdb;&=SX1QL6G]]=US(MN4=RAIYM3F8?+Wf(P=>+/+P2F,.5#VG;/AEd
.N)1a7LPHf7ObOVB6BH.Rf2^YWP-KE4Q[1>)a/RYM8OOF02/-LIT_,7^TKa+:0OI
cb5ZR#eZ:KD6@013LFDWCO0=;(K+K=MO_BBT#e3f)89^BVD8P1DN6;)F7CKHRSaS
9>>^MRc,O.D<Ic:.AFGB,S?JXfD:OcME(,H3M3c8&ff>C#J\^PF4PC3,d#[I=3A^
Y(H\O_0LNL(CW_]#?HC-.>RL<C25I=01S_>J?B=.W3bW(Yg4HI>0VB(-R7T<7YRH
.TRQBI6@+gb.O_+W3Zf>[#\e\U1aJe/M(eb<SY7cZ8&^M#X8E9VZT_Y,Q4]SHd2U
41ISZ=BM50>7OY7BK6/D>c&V#T?gK_QV-/,e43cGXf6:>9<[W32;3#IWF>P=1J_<
,^6BQ38PXfaaJ3fGg5S;W;+FCXf:Y8N@3N)HGFU=.7b<OPI\6.37YO_)gBYC2(Y]
D=Ze:A2:P<fY@e\37P9JS/<=N>5KU<JNOZ-Z?,BfC(U5H4)eS<Ye#QC)RgQ)53E(
M>[VUDG?fF\RSa&07SM6-J528B5GUJ(J0^XWP=?8NGK9)717=GQ9PIAC+;d9>0eL
?eZ:dWZ;1aFSMaV#+8O>A+e#H;-&W_(&0aGRQ<>VG+SC?(0/[</2dL3?X/WJQ,9^
.<X_^g/63DU#&Y4=/Z<_&<[E=-R;+0UM+.>\b_SWY[3\5L5\(TNgSH1_;bNHCR7>
WG;-3NdP^dA8X6(?<V;Z^7(]5SP^L4d3_G([I];MIXU]DJS:?ZAM1.@d+7]f==5N
[,.<4P#,6F:3Z^&PQ=\W>_S?KA]^Q\?&Fg+WWY.N8Jf;9HBYQC03&K<^LUK.ORC8
SK24d9d=fdg_316F\cMBZOad^McOO)M6(:I[F+YF3+59\@PQS8M,VOHcPY9U8(5/
:7R=WXH.-Y3&:eIH2fT0D]8PH6B4K;C@Wgf\g@g87X#QI.6FTJ^-WF[ML#V0YSeA
d:d_98)#XYRA2EQ3_2AU/bf;=[</Jab#Q?91=O0=5b-1_^c1YDEFD?cFO+C:]RCQ
U9H8A8-Z&(VZA<-N0L./F0UYLN3B\XMbeUVHa6KXQc^323J;TdI@0X<9@Pc_cSL2
4C>bJdB=eJ=4D]<56:GYg<BR&+A.<Q3MH]H<O,:c;;MMOI4.>b)4PA4]4IUQNK>6
.SXd?;;Z@LD?L5]PUaG9VB+<.-]/g[^e(#9O/>aMCb5EJP;^dXdGe,:Id16X3LEU
V5Q,=-cK?^INf\HVgEPVT9=U5983=cc,Sf4-)#&f6BBEA+(38&4<U&cf@54c8C#T
_RVVM9fdCf-<]4J,L0G\3HJ3N]Ib2>41L4YT@b73-Lf@<^4cJa=aN;+I^^-.g\EO
g=BVL256CTU()9RJ#M3,aXJLBR6RD.JC:.QAE,>SJ?<ZO4-O6D-T+GDRgO02.0)&
gIKH>-c/T=\CGVbXH19cDAW>?P\3IEa3\U)X=9:/^Q<90F6:,c]>DaCMb2>0H3P9
L=C&Z>fX.Q(e++M?N+SP[BMgg3R><3G&2#Z:d3^a3=H,SWX?96IF>Y\7Y4R>)fR5
@\O)Feg,+=eNT0NX/1XcZO(fWLP4G_MF];Z9TBd<Yc^7#GQPeBGTKP#K5U8:K1PG
#YT7MP7/5a.<\dd_fc2IfJfJFVE_O:D>4ZU_KbBR4=/KCE=+c[1<e8_XMVEb(g:8
d(a7RE0&c;T,ZX4EEg_4I0c]9<H0-)SJc/[=2=D0NS]a#6f@:IKR5Bd35YY/_ATd
&[;>9REZ9Ca>[]:M9@?7S(]aYS@>f?KG):,W+A8\6VF>K#YRPE]=O>N&;H6((AU3
\7XM0/dXA4Hff^YCQ>,F(DReAC=(JT3ZaNF=9G3=O>D5R]-J>)P9Qd_-JaYc1F?d
fC9G/RJ05XI&CE62SA7gb3VYc;U7Lf1.gcS1ZAU06CDDfLWQP,#?GO0;OdY49<-1
)]H&c2<W6GR<5?F+4U3?WW;)7Cfc.Bd<9;Z1X9:bWe.I35aF3L/.9/.Le/(O4.dK
GfA1\eJ^dT?\/,+R2YGE]e8+777>HEd#0(d5Ve6=41OJFXPgUeXPGdET#9Je\KKd
V\F11755@GD>BgM/U0cgI&4/OK[]IDA-VF-Y;M6K3TG..=TB4YNNA)JJN6LF\gEE
&G6aTc;I:4WY9)5T?^Hg@7H_ga:e.3X;,5HW1?&2DK[:WB)K78Af<5.6_B;[QcA.
<,QYH(819^+\]\,V7J@VA-YC@/a3BUYP5+cf_e9K.)(0^1KbW2F5e43>bQK.E26>
H4@#U+HRFZU#_^2.-@a#([d6N&//ZM\e+/GKc/1RR)Ae4U&Y6e\=dY<S3YESMBKS
=DZ\PSU)Q0bU+c&I:B18-1Yf?8b/9TBZBaP[LMJW,1\)I<-B8Bf/WWX]]g2e[)/F
JIMe<&4#ZKXGE4VBP\Za<:A78NTg;N&X3Rd?CT/TCc#A2AHMJ>&=,ILN#R22IAeK
XG,E=^?OLAWcO4@;D5-N6g:1J1EQGb2Od4SMLV]Tc5f-/113,@RB/5R\DN,Y8=b2
VT#?MJB;>TKK)_9gbd[a&ULL[<@7:1GHY@\Y0SfW[2:6DXZ#GWLTcCI,=QWbCQb6
Z&TTCbG(8>BOb(<-@cS4P<J3:,8a>P:7Q_aMUaGVd]#Z:MbePf+EVD5,Q/7TD:Y>
WNg.Kd46Id3AC3bH>F7e+N;E+B::;E&CT2V_U]=Cd+/[5PePa\_@893MDB4&_P^F
Fa970.D/H>B-MUYSFC8S^I<HN3Z\bS<R]=30=GW<@>T:WM\RNN6=7?V@;ER=-ZWb
_7<AJ-4A)&a?0af>f?<R@QHbI6[++#gYf9Y;L,4\[,N(K,bC5b:;&J]H5\2R&0@>
\#_5@&/8#EWD:4AAF0eO5R[Wf+\<aG#Y>6ZCZJ9^S3&eC>0Sa9J[6MBH+4>eU3J8
SI+.JOK53g@\f:<B/:F[VLCg)@U1#3@_[8+&.gB-IKXW^1LO#9g]eL4WTR7N\dVO
1N4^X(8Z&8H-W+afQ4-=AR?)eV_dg8R:O-2\a)dM)c2I8Z03WJaS)YZ8^:J35ODN
fKMCYb)SaR7]dbMBb)_fTU]-.7QXCWCQ;46SR<RbIENSZ6@3\NZJIA60[U]gY/:^
Q.#PATL^&+]fSQ9Ud83Gb?C#</Ae7baY-a2&R)[\IG-(&ced;@(Kf,P7#B,+(&.@
U9G@fSXJ^S&,2gP9WcTXFU4<]Y\0OJ6Z=C2:Af^;K4Z8T_XV5IScg4g&+7]FKIDE
=8#)-:,T&D#0Z))(5]e-Y6EMgGH\MXYF6aW@Y-+ECBESP_>^\gQY)H^PFGFZU/>f
CeY>E73_c?Ybb&44fTf?VP6BJ/>R+6a5;2?_Y;WI7#+5FS5O+-Gc:X?BF17MGB&a
&<-M)-<d[d?R&P02=cM^T9ZWaSb;B_DB,I5Z=aXSJfaB,5]L_dKgKe1.A>WQ8G3b
2I7acBc>Y@D4U>]c,+R&S]aM6B1^U2^cd@XeDd1@1Bb)?K@<SNCXW@\OXb1/K8+3
G85-0f4a9QJ1Y6\/04V.7@SVaJ],:[+JX0GaRG(PR&Z]S3We_R]ac:&]ZS,F\aB,
55WL_W7:&;0X5)Ogd\KEdV^SC=K_8@ICV3NNQY(7B-CL<,GUZg-(c_7GI.X6F;@Q
Nd87SJ^JDdNJNS6@]=e(AJR?A>;Y+CVC5_KDORV#15RIB(J]H75FNV/VcPSC]4Xc
?JD.4&1&V]gJc.S7I@^AfC@>_1^TV<#dCTG._?P01Xc(]&W(:g9M5.^V/J]6Z::.
[NHMfKU:1XTA\4#Gf/R5;7PcU4DHXY75>.INIA0DU:a=1&+O?>aUYK@A4S+\\:\^
=QZTUS6XeNKBO<5\8,@KZMONHTW?:)@HZ;S2S#aI[Z#@5A0>K2K0^X1P)N.PE2fE
>DU(4P@^20]NV)RHaC]g+QCLc..>gW#cVQgdTIb7Y8EMYXDM5,(5<U9G(E=D[EBD
;[9L)Uf5O:X2_a4Md7>:[780AT:8,aZ@.Q>M]a[16WRN[<9CYF.7283&Y=FF5XV@
.2I>>RP1eT64V\)VTI/dENM_V1UfBTSHbW,9PX2SP:HdH:_QX#.:J]KS&T0A/^2A
>>ZVf7HX/EUL&UN[,_8#AfL[PH4gF9A>K,(@eNT9<PACV^cfad586SIY6P6Aa0Pg
(VNLF9+g7aC?4P/4KRe(^[PXI[L.>Ncd8.]S6JbX&OFLW<QV#BVS3PI)ZJKAf6:a
@Y+)1>-8OR6BRgUM>\e8H?:WbA>A:Pac@HMQ<8HV,^-LS]0@0W:Cg)O#[DR?@O(0
FG/Xg&V9Z@11<^bQ-^d71R.Q?,Pc:C5]fB=;.(KEDWb>6;K:]3MH#MgJ[RR0]6DH
;U2\XW(gV\g,_EdBS:TLOZ2HE;\:&ZYZ+4Ie]GN@3]dddH#CDAL_Q1;;;6:SNN+5
+E->:X/XPPJ_T1]<>NdZRKac^E,HTc5-9)fWd+O]K,6:;IZ1_Z7f63IB[B>6L/&H
-aWKCM=:U47?.>SK/7+?a[HHIF+]G-,N20?62-N1Y;gafJ(PZ&Y@6QO?DD]A>ERD
[-W)+Ua):\Q1JIU.f>_:SHaR3]D3Ve8LQ3UXOR_U2F6B+UXfUK\10YTeZ&YdT6FV
E:>PL2PB\1>6g8SR@Q>E?>>.Z,Y12&&SFfJ1_\f8E#PI#?9DE,fNDD^8Jf3P&Lce
G<E&>FL&Vg,P.3;M.WV&99UU]H;<?-:G4<JcF1WYEX/AJ[5QES,b#_6ODJ]YbQ/e
]CGV)[-D3CDJf+3g<E#:@W>6H<,6(&#EQ5H8JY?_#e+-YL.I(VL/:^9(2FL)(0SI
63&T4I4DHCH+)AU<0d<C>E2VC&5b3cBO<8RE:NKY6G@3,BS6dZ&C_QU@(U5,Y)]U
U5Fc:aWGQ][,SOTH:@V#99HAbPU4/G/S>bBOCYYT:X[0JSgLa5S9e1&^MABWf>Q1
ML&G3\LF]Z?>WE45J_Kd&G@e68ZIY:+6#NVcEP:P9/060PZPWU-U@;E6]VJ7]Cb1
<b2g8,@,7<9<JSX&7;_A]QJc11.ePLXF/N\C7WWYRFN6a+3,@Qbd\1G8WDPK?LON
C4SV9JOO:0B642L.Z\Ne4SMJ.5dF,.\3H6(>CW>QE,b?(#YD_=H.d+(?ZK4g<,PN
8=eg^JZOL]JY/9#:bF=()7,M#=50NJgY?2D1K[SO5bDF-/g][HFR#67I]J>1_JOW
9(^\W?NS7TP+OWT3>MN,+>3fQM?+KT<O_PTc#daXG1bSgAU:F?DZ.>FKZ>R69QMK
,f&9K7L2NNV->c][+;:_BM#^B5XX+,Y>&JC4OW#R8)YK,cL:H00L3MA=;XE],9V&
HC/V;IS2Uc[ZU[+,5fKW<P&CgG-fSH>(N]Z4@B/=4[^\7Jg5Y\@:KJdGX1J..aaX
<TT@aHK^/cc2N6)]aQKAPMSJ-@X[>^&Ba+RdK;T?ZHda3DVa9F=,Q>H^.PFWa:W2
]OBGKTg&5-[?]VQQ4P8^JI#0XSI[GK]_56?WLK0U8c>F5T+(7T)IcJ;8V+a82H.\
99&9dU4I?G11W6#1bW(-g,46=ZPJPag5a#6#^ZC>2(f6]4MPPeKSAVGU?cMHCG:B
0e:,7IL6-Y5JG2Y4cb-C;aB6W3]JUOH[f@RBg32TcU+U+C?=PYI[L3c6.#ODfdB-
-FA886@WA(:#GBAS1HR7<:IN2RG9ZO=)#1;(>A?)>;>@#Q:2IAH3eGG+Z(:WVP#G
E&M.QER7EIQSLTU]NO?fI9,YBT=F23>-HI5\QdOQV<=E)>QP:cS.ZUb#f8Z[-3:X
3NLQO<XS:IGP5M^R+=Na0>R70VW+8&E26+#:][:35Lb]-MNa=AK95eP=f8[/FNL@
1<A>:Zg4:]&R<YT?+,a#<1K1_9=7R,eaI:S)XR57?=a4)=eP=eb[J5g.BG8Ga-E4
X)?]::cZGX)&;L/]g_?VXK9O)9W#XOZEL(;/N4_:_^FRc7JXCN+5Q:),dE-,:J>#
EVKRC.NJ<#9VCNBa#b?IVJY-@2_+9M(Y;R7>3aA&7WS-CP#I0,&^/JANUD\HKS.Z
F3]^[BOVLePN95+&W)F-Jb_J/?IX>Wec[^P9>:9_1F1W27:4H#W#Q@7-/Z/Q-MXF
)Pc/:[dTJ^bATO<5[#;WSQ.T#T?+&8[N5DgWK3gV+_+K3)#&X(?W\0Y/H,49Q<8P
Z_22\86QJRDY>K\@Rb-VgM5DHa=,>_/dYB5H=[Z[WIW85,5<Z(?]W-)CUa6L1?G\
_BDVPFDdg;e?5A8KW2\]KFV\MO64JDPLS.7C,AN&cZW]SX\KVF:1=>S[N]U4cYf:
-9.H=(2_HL]g(^1]4@7cIH99-O\L.7IKfbA:Z)c(\X?Y,@VO&?c(/1/PKP.I#TPe
+Ifd[(K)Xc5D1C:Z7?G/f?WfPH(23Z:,O=137<-fLd486cCM27?)3H[5d.H\^UN,
J+B4;C23KCF@;Wf[K[=]BQg)41O4#Q^D/WNRUHWXY0_U3B];[#^UOC=<TcA(g08/
g@VSTXCOQ,PH5<A07:8PdZ2#PK_0P_7,NB9>7NESW>3FPARWgaY^Y:\^4\&aXSaD
6_=^-^fB1E]T8@8.gXCPDB_#.O:aZZgg]gJKYKW53M(c&A@[[NIdXXP+-^.J7eY)
f^MG@Df.\:R,+?\/E5@2>3I^H97.2O7O@EGXZ:+H&f<8ScI.6Bb)bV4Id)G(c#_^
9OcV&VPNL+>a]==Ge#R/@5^8WRB6[3L^S+FcG@DK3B<[4:Z(4)/YI=]FJ&6=#[ID
(.dfA]88Q.(ZCM.I)LgFbD_R\CJS+dZ?Z/XJ41/2X#[KH1BE,KSJ[[S6Ze&Bc_]&
]]QTL>XFC0A0G><7bK=OfcZ,#Z^cMC5Y5U]Wd:d?\eWCfa+^(GSD4;GGX7C85@[&
G[[(E;ZMNUO+^U&4@5AbLGW(]<4)VU]TcS^<EbO9STZ7L7d4?g8<X;?cB#K1E2D4
cOgYY7M.;J\?O6G0gCC[bQP]cdJ[,.[:UCD,_gQ4INS+UL&VW<VJ4E<U_G>ZZ)D9
S=):W:W(4Pf5?D1E\<N7WC3P,g6K/UIbK(Uc6g&>:a./7=[YZKG(#S?;&9GY=]a4
7#aRHe9AbR1R^MAM:Y>gPSPR?/H_W42:P0QP^][V/Q1-FG8+d^=QJ^1>agGDVLe=
H5K65]NeSc8ccCANYAgAZ[LT&QNbR_08VAT_U/:3L/1.aU;NF-PK?cGGaBR3>1RQ
0[8\b/Q+P,TS@3ABH,d6WD&,g<9>6[T153,1D,TRaaeg1,cbA;fVc\bEDOY<J#2d
(.AeGN#g;AZ@E:c+0KHcY\HN(H9BJZG:J:D0T2OZ&JeR;-Ucb+R^_JF3/;SdYXN4
U9)Z&)FW9:W3c@M;?DKVRV[O<>ON\^&6c6)XN?fOc2(X;B.4A<59DV#&>TSId^5[
4>=H_7,C7]b6U.-f>JK09VaWTR,<PPMce)/3Z&H8B0;eVX3.]TA(#T)-1:@IT&-:
_dV-JTQJEVV#OUf=3HfMBT&1RV@?HFe\L7WM[d30bAHXg\2Z#0TTg2JJPH.dca@Z
Q2S8KGg]2)+:,(.K+Q[41YC[ZZ4ZL@UU.CT05:^^QfE;b=^#Pf4QcfTg&gcXL-5D
#fF\+[IN@P3@D2a<HSJ+g18aRZdMA9A+FDBWAUd)2WFYSg2Z<a&@5^,442FeU<3,
/6G94Xf@@?YZ:C&#RPPQX=KBg@[]X-WWAF>-DNPUL2IeUM7P3cB(R.:/X>?^->^L
WeBP9,Q^.ZJ8VDC./>BRffSAC6+W#F73d8UX9R71@;1QYee,NUc=;9Y+7M9G=RLI
aI\>_RR8H0XD7Y5CMQI(\OS?PLIN?dV(_\N,A=..BWD_,3ZGE/g=253JUFg<G+];
F0H>g7dJ>;)GO+-0,af1NIGE?S5&-)FT.7#)M&X2BL+&N>^;SZMYcAJ&(KMTW(^X
J(aRbPV\EYK-QGa8eL9B/b#=#Q^#X;D5N5g2U&@MS;Z?eNPK3,3E8N1@d5QAB.fU
6-US=W40W>cN#?-]K/,d:f3;I)5>[@QLP=C9VB649FH6I#S,]._-d9KH1Pg[87e0
1UN85^gM4SDgGM)6SF,>2AeV8.YgH3(fHHLR56Y5S<bH+S91eEY+IEBB+ROHCIdT
DOb#-Q#^dgF?:>?5d1:8F76)R2DcL:?6NC5;.d4SeIRV(aH4H2D0=a73_K-XU-8L
Gfg9/,7NQ+5YXfGg3+Z+C;[J[X-@De@^Nd&WVSEG-K:C5O17A-#@g:1G:SB@@,-W
SB7C1&R&dg4)/W,)OBbUY:KGK@FT.,7+V./N-W9Tdg>d>23@c.?VW-QKIQ.//WJ.
cgYOS]AgK6GEd[B_eB#QR9.V/EJSDLT&GM[6^8)e\@bB\3MX]bD=P@(IHf][BTYK
&<TU9,VKHQ2W[T?gA/fT(C:A=-85f(ER;,gg)J)(=BS6M^A7+HXX80gQ&I<6RcK,
bH2T=0QYTeO;3e/S2X&YD27X,O^)7SE0ZP:SO+eX6b(fP(I/<TUb)e#JIR,ETQ&D
S:f5C8]H]7,PRTTd,JIFX;MCKTV/^R13B(ZW1.=G/dN;O?bH&G+)X#>?WXOf1->9
^T2MLJ(UNLZ90?&+;L17H>cG&d=QMLd6ae49U8Ia\SXc@E(?WIc1TZYJK+?-SZ3J
FOA+CTQa]K8&EcPY5[)SXQcP/cD_CFbE10(f>Xc6H.)TSId79W?OP,A&fP396W74
X<PTHa6V=Z6BV(J,Ua0cD-D4+(GV15\F^E;55V;b\S3bbODXM8F5B6[WX?B9A-5Y
LS^-X5@NLF(]bBSFFA)WNU@Qe>C4IOaC&,fYU.6FeA1U^Vf,2FW2NQHeX&c9@BHB
4d4Q\JZM8[FLU66-/WRbXS]YaS=)8c8>AIU9@+C[G8dK-G)+RS2S+B764g=2B&Zd
MG0#9)L_agTLW2#@0T#W7cB5Y992/b(cE<dT^cRPZ)7]D;&U6E/bgH0=.<d1U-g9
)[N.-c4[F,bGC14XQ=(>(@4g]g9;]aQIJSD<bfS+_BB;H)@)A-IY\243XcVa.RG2
P\J=SaX,NSB@MAD^<9;.OJ[NeS#02H/X1R=Q9c7HI;)dS_J?b)7Qa=T_B+3a1e9D
=/\[\.26bH9G30UcZH5V;L&#b@W2T,J;cIY),29W-@V0>N&gTXYFUH,94B2X8b[,
WQ?(\-_ZE;(<EZ-/15&<DH,\g8cAL#)_:Jc#J197LHE0N?@DRcI[A@#3ZZJK63BY
I3>3K&]U3fSZ^cU@C4IC783DaIN[/\3MHg2Vb:g,gXXEUYKBXXW<4Q3QSL4P_>(5
4(-5\AWW<:O-/R,KK[]ZK0_JZ7gDIB/2LP2(KI6JW5J,VVL8<CPPf,<<^\9O/<-I
H0T;AS>#2;_V-ZR6N[a;6[4R,)9WGdIDN=5.Ig8OR_]?I:dLJ0:eeP\&LKRAI[(.
>.0A+E@0#7K80:AFea3)7L.;K>D0J<:^S_cPDTOQK_eFJ#\NF?</)KPK2[0;_L&F
:f.F29Ka<6/2W&dWG23II(/9VZ\4Z;BZKI^<aM\Qge/JZ?HY3&S278;W?/dA_aHK
7:MSB+#L7^A0c;-:.DcARJ)9c0c.>0//,+PbW^GP2_1Vdc19,1N@H?Z_?]8DXM7:
[&(^I2V5>W?Sd@CRZadg>5BG8cC:Uf+J5UVcfH&#GA+7Fe@abK+8<c^E4=F-[F)?
MYfT#5.K8:2)?J0PgOdLa(deY-D[#=],AU/,E@([AcbRDbUH.Kc^\\.<aO,ABG:6
^T(?gR9BOEE<LV)Scg2-X2R^<8(6V@][Ja/U[D#.L&X,]MB729KPBJ1G/Mg?,b6g
LPMQ;f^X6RI\)K;;BGe;UFJ<FfXEJWCRBee^O&cJGHE2?QI+g,#-0J0)Z&Z[\;DK
^YcEFd1Z7/KTSTb,62E+YZ7bU;cgF[b?+(a_C5@fUb._>e65K_^f5ObI&7aIKYaa
4EMggFGJ==4T,QBeC[()302P=@GU4W4&;VQQIVZe3^=6W9XM&[ES7Jf8EN\aFQg.
Xgg]]AKHL(OaC/GC7^eIM=#OGcE6:O?HE:&a91?EJG(=AU;?5cUdRN3\,WU/(B3I
Jg<,gV>DdT6KZ8B>U4\@YU=C=W4<a8_6E;&Y@O?8gBJb#HcH>X1M.EDH^[RS]<)&
eI63979I1bG\1DHS8e\6S<G2MM&G@f:(F<UQXA8U&(Z<92LB#34)QSTFA?(C0]<R
AT(;S<S@:[=]+W1:YG(<Z#(6W2TY3e@&<[CRQ772J6+fRIX_ZL1@&+R9X96]J+,?
B9eU:Regfb?.DSb.Pa1ZDc;a1b;c>/aR77>Ude_/87N=e=bR#aM)JO+G_M\NNNK>
R7^E&YVZWc,7;^bM1gFRGT01&8c(0V15\)]J/4FH3U.[&TNL>EG2=D+,9Ga:JJd9
;L.\-H.YMgT,&OE\TMD_.(.Mc;ZGLFHXR=X/aB&96<:D7H23EG^@&KeY4MK<a@?1
(/RHZ.:Y,?JC0)=N2)VeK8B4b66IfL]V8A2_S[>5I?/I1Xe=4OQH0R+QLV[MaI?^
&DOPMT^#)31=H9+8KNFA-;-7a0@M-7BN7I+QV[C)UY^G_g._N45W(MN(P[O3,Cf[
6>g[D497DE2:d86H)I30KE?6^GWTVPA@8,;W>21R7XM/,XJ/MDO[_@;&>W/1]X6+
-@R+FU>LZA^T/aQ)eRFYGB(/=:U#-V(2+8:e;3RFY.ZAL^CH_@PcP8JCa)K&SD]X
?N/&I^2OXdW8M<MR.Vg[SK<J9F.dZ#UOQ,H.;W>geR=Z1@MWZf&d4M@c/-ECCA\a
-Gg;;(Ia&WB+L:H3G&V1K3^U=J@H9P[7U9-2=]T[-e[,R4<9gK4I@Gc(0SfSb6C2
eJV^6E4Z+Q:70]MX>HY_@MX><TW?&dGRS?=E55Z#&/f0,c8/W,Fg4<Sf_C08Z;gW
-8Gd(dTcB]\LGBUaN]&OJWcN8./OVPb-2669D\XAEXBF\&;;>[X[[SU&LFb4:S#J
__Re2DeW&?(N,IW^>)YA2R84cDLBW5a.U-OL&gbe?WH#VGU5>&X5T?NS>XL1:L;N
>Va(,V<PXN::1dR3O09Z_MCBW;1&P;F4YaNX6IJDYeb]<_)f]ec1_>c#^P>@F<QV
[Xb3,?61E&;K?N258-_gW.5MN]+:Q,B]V;R/TEKFFb\a@UUW66IW6K+_HS04\T3M
>TG[-1aRSSeNIg_75LBCLHBeI]_U8c7XP#:<LDd9DNe>B,aKKL2S_G.8=5OQL.C4
g;a[b<UX\G4VLIWZe[f>3N#Y:T3UH,eQcU1HRd7W@+dXIG\VEcXDY5fDHKY4&E/N
#X0AMb^NZ40O,LC66(J,=C-UD)V1D&KZ?Xb;+J5PI>/Q>^-DYc[\DP^7F[3-d(24
+V1<C)d(S9B)KCL@K@:N=V2,cAL.dc1MRgZ^8EL??5)02AT3[)VO9)PbM>da[H,Z
+FDZ+-[;;PRF+#TOJ#<&@9=^GHa_?=>P>@H-563P_-.fS#fSg/=fN2bT7[[8I4M.
L2H&<,_Y93#0?G\YgF#O9SdK]R]9E9#KRab^f-[F:#]De5^SK(A/0E)85-GF(WNR
#Z-:,^bX/_VBZ.QV#H)Sd.5IUL/Q\5/G]:DP\,Y5Hb;f1g0cVG59DN-@F59S&1b\
+,[\,-O10]GTOb\B-=d.?d/M(?\^/K;OK&bS(ST[D;QMO+(T=7O_Ie/0YM3CT2Kg
3P0+/A=NN6QH14]/_:61M_I&fT3g=GU+/=93df&Z@GMC5@3GAU7\\[K\PFIPSM7,
.IcE&8R52LcRH6g_&WRa2+:[>-[:0\<6bf30Oc,=Wc2[d.)0(VNX0:e(d<dVTDNa
?,_#.;AKeX2YgN5M;+I@2A6_JTA7#8@U^e^UC9gG28bWZ4Y+(Mb&WC=cI_10TQ01
JI;QD2cJbb??g6;^&70Q#5XNab:)CPLc#[[C35HbKPKdGf/8\+E^Ug2RUP:[cO_#
&<H-[SFDN_D(P6gg(Hb@ba9WG&<K(=)VOdD?cd-(Y).;1c)X<=A?f?Z1gX,\>M8L
@NM;))faAQHe4EM+SS80bV;6F1],[@40I))PVX>(P46EdZDPBO+19<+I.-f9,H^&
K4N.T&dM+&[3gP5D1C9gZ,_[=P5:&_=Z79N?HJ\VK3>K1ZE+^]UKZ:He6bS#MF+M
fVFU2:Z?^f&&FE@V,CG0XWB0?)_IB&/[UDGeSE5J<8/V1<X;I^78/;H-S32C(6CM
)I^_HUQA70cFE&Ff])+AVW9&LD<QVdT-P0[c+/:OR&g4]G,CW,(_N(=\T.QEAc.a
5fR8=_aPZ/G9=;Z(GR0,4I7N6Y]L-Z>Zd#ER19L4,-5(F(U4);b,UW\&U&T;@g3E
=ZcKONW;QL#H-)fc:Q2MW8JgaMHZ-X_45FJ1R-1U=-3<^?P&3_.B\_H@TTABdUEW
JG5N,HUPZ/&ALe&Q=X:WgR7IK5VEH0c=g?9?I\GL3D^3:L+_-,]9RKR_Y[LdD9L,
-LY7d.6He2ZO>]?g;EF?,>W:1:-BeYBd+AF>6)FTCc3bE<69Y2OBeNK1QR66WUG]
UgQ\:[8/L@OcS>2\EfB-KDb]](@5+Y(9/^cUMSS@Y>M,E6,J[d@?61H@8F>H,L@H
OP,bR6b)e6>\4a9[K./S8-+.0:#4#,DTKU?ULOa#>M>;23Y74[.g&Q6C/CDJX;XR
Hd;5:@L0?Y[e/7ZU8KNP+90O3BbI72U>&WR#E5>HWBcfO\6DZ#e:MbX4VU@2L);;
QY=C3FSI\A&_=,Sae]USJ95G?2AVf0UK&;M+Va\d-SJI[C<PgQ3@J0G;;/6CHD,G
8#02L)D[F@OZ6,Z]MM:M&4A8]=K>WD_;-3-?2QFLOSd0A[-MfU7J0_INg0a>[3Be
3X]d6O^<gX?/-VHL>,a&<a?/+fP,=)PX)E0N/MVaeHZdOAE/Y.L/81&0?@R_5@N3
^Q+QbMV3YaZ/.ZQ(aH8PeG#F=)EGUfH-Fd@8b3>=b=9B_E3(T8XILd>,)ABA\T#1
=NVF6QYQ=HDYU_19:e)7-_Y13B5P(c.R;Qa.,A+W3c&:1X@@J8#cVFfUF&>0PcG1
:OegdP/cFIaDf6J/d]g:\a[H_7E:GMf>KRK:130B:.@220&_9N413CPc_7@5[UP5
47W_fP1a\Abd-P[#[?VY(d&OK\6_>Rc1SB(+U2f^E2&L;0V67[1,M\KKO]3e6MVa
Z,GCfXHVJZ4?MZGHaUET(&RIf56#T5GZYU]_]@cHUZ_a=Z0S3.#CC9cJY+Cb5G]O
]LGT&N8R/Z++&QdgR[C#0S?:YUeb-?1@W,@bS=+C8V[7[B1.AN.&<77W:@OQ#81[
VVeI88(VJ1BC(E=DO31?]?_TOFDL)]PgaM+_&.6YPSPT#23]FcGTWaG[cI@/ZE:b
FSE5.N8RJc@TR4f11C<Hd=#8#?U3)U78g)DCT@IK;FbLHa.Z,W>9;+>QBBc+9O[K
fXg77_=.?#B..D0S^(=?H2J-PfNae^2)P->HXE?g+,/c@]5fM940@aNBSHb]gSYf
DLgNc5I4.^HDEC8V?#BG,A1MaA.XUQKWd5fBIFN>FSBS>e&d8]P_\0R6F7^Fa9L-
IAZ_.L&R_fFaa)O4P.V?,aeBfXY2Cb#00U\10ZV;5/JYEb4,?K:XP^a4c.cgCF;G
5#E,+2O^FV_D)Q[.-/Ua@V6LP_ABB9&L4RCAZ/5aD3ffQ]EZ2U;dUU7:I&D#<==C
G/XAbb\d&LJXa2EI)2+?V[ULIWQIL]X46X3eBgUJ#<dY)_K]-162AIPKd.PT8?eG
]>EbFA2OC4<5R[/HWJ508\[3PXG9R;<d+2G)^DI[g1KgL8Y:6++:<I.(fZ6I^b/]
M6PY>P@B40@2/.O9@+F(5e5-b53^(8-WKYSAX-0R<6A/FV/E/N#d:KG^cNOPG/BQ
;>)IN&0KUO&d+H\YAEeM(2(#V+N([d\e0U+L>8<(I8Y=+GO/U77-:(^_VZgXRA9]
+CKb7JZW7.C87Hab[3KG)a)Ba-1<??B5^eaPgc5gA9ZK>GXY:.e4;UA,LQ+c>.WM
\aGIBU=E8c/S-H,I.Y6ON&LB^;H/e)GbUg=,EE2?H]W8PM_;eY#.+2E6PDfBJ0<d
b4#HPeG>eHK59eBEA/XZT#<)gZ69Q(##d>f9@3fA_-4LEBS^:=:J)9@<:)4R<&4H
d4S/HO#7A_I(\N(Vb6;<UE3IbfcQ=d9V\VFGUUKV)7c=RW;E28P(e9-3.-\EgU4_
>V9_.:0#7@FK>Q4N6TO_;MJ.N_]Z3aIGfE.W:\):NF+UYY-W^Q615c@3,#d<01[S
3fYb2U4.>_X3b(c6S2OE4^ggRU]AM+-.-,CM6b=G;d7ZFIfX^H;8H/+\7=Y;@LOR
F4I]@fL+d1VYMW6&aRAFQd,19#f&^STCA3)50+4_EaU6Ra-U\6#BOe,Y]?/8-C#.
Q1CROD)R-5W7X6N_b=GOKM4I:/T?&.JAc.Q.^7+UgI];FS;<:#eb+&d:b8YcI-X+
F^(OTPSJ(bDF1a::&/Q#9F)Y2]Gg??gC+NBdNDFPgMS>Cdb(/Ze4,WcQFBa25J<3
AKYAOD_M6?B[Y5N(+LXg+UJ25AHA1-.MQ9-?>VDc[DC&K@LKM+7PPNV23_:d35^X
\-_aNO/V&YH8e9@0Cd8[2IJ-5eSYYNeag,IY6aKEL_=gZLIV#/P16<(]N@gX&)(B
QF:9)];UXW8O0VK/[YY0YfA+VDV(b/JfHI=eZ>=.1+HBK-Q1OH1[NIE=J-N>D#/\
G6]Q8(J5XF1(g?Ce(_6+0[[W(IGLHJX>^EI?d]:g=1-gAX]GcJ-96./_X;GI@9\N
_H]7PQ(?_<49S-N+H:H9W/gDgGf>I1F9R@8OQH,?M^RH?\Qb0?V(BDGTWgL?PP@F
DYOLRBD(TKE_RCAJ1Vc,HZcgMQR@QTOb-df(B7:R@FG-1/JZJ41aC&^f)gWGRQWH
a>>/b&/D_H#ZQa2e;G42)/TbB9,EE]BNHd,+SLJ6E@;<8b8HTa=Y_UcC89V<A@Q9
(DP8P-Y-,I[/=>LYA4QCSRGdgUT0]\#+dL#[gO88I;V/0+FaU7KE:0?X2M,\WO2B
46dX(7;ZLc.39.SU4C8<&B&3a.;-[)YC<7fdLG4H1A50@BKL2Xe\GJ)2-Md.M3NV
OY4Z4B4:V(1#NNS\#):NW5aWd228C#,N,RW-Ga/#)_EeC?Me)8X=>VW?H6aZ^Mfa
>f4D#\M[e7-/C3OWU@&;X@aDXcYEKU(a)6Pc4]&CN(KSedO>Z4A5PL-)QU8\H#b3
CA<[P@+_ZPVE3+dTO@+2D[@YO+M+]D>X48F>7U:&FZTa@a5A(ZgV^7=UAM^bCD8N
H9NL9d\+4-d>NSMOg><;38;-G4911EZ)]/+d(d/G;41Md7c^45;3c-=RU[G]1_?:
N7K_>KOZ8+a4DeT4,;:5JX[De@N0MBKU_XEg\b8&M@9?#OBf+\KY]7cG]DE84E)&
>J64g]AS)b#XdJW_A9[]=^AD>35V#7^>:V_f7.YI+HLc0gR>55,6CD27WY++cIR_
gdYMC5K\d+&I5(AgK>eV;T\b1-GMEHTG7TW-1bH?1,<1AYITM#FM]8&Q&@ITQS[d
YJ=20(>OgfcRRDVA@\\;W<2cT]>0CGP3?UK^@LVe<dTVA:-41UHZ;=)BC:e@EcWF
8&SD_BT1#(45.P5G1S.I>HHC2VbX(Z(.Y=&]WA[+B[:L75:a4PTH/:=PF3E]QO7?
SbO.MbY&6Ege26Ag_1I2VVc.AQ+_[XKZ5Y4Y;NAFbXFY.Uc=8f63UC6IFNS9X5G:
/0/aR[PS28D7->O3?:[gTD[cb:5^47X(?P9B/78AC[g<]0956E0HgfbL_ZD>+O]3
O_(@LQVM>D-I1SL?->Sa6KMF_eAM/gK9IN^>8NKN6Q-YGW3[RKNUO:WELfEf#9ED
3+J(5GQc-f5+7&0?D@P\O4&b/]1U6IE[<&/F00SD15b5,95ES<6_X()H5V6>3bE_
=0<V:260S2X0Qd/\H>3O):5E8F^a]MPTZ5VI?>HWJ5?F/22KMNW)D#:+HYF@5\9V
6)f4M=d5D=M79@_BZUA?ZB6MWH\AS\6)EE[#e&>W8_Dgg_-R<W>/N1=6I62,B+V>
e<^AUX9BD20OA[T?@TTB-g#T]bLCfW0a_F=HX^<3fQ>#5@16GJH-T_WK8([X-Z2@
84QX;XIE8,?EMTNg;2P#\R-585<9P9g,(P,I&O2BR4.@?=>7#<0Z;fAP&M/BHVI.
LEJ^g+SZ6VS/>OMGZ<&GOQKNB?,<eA2;g&^Z6O@Zc?+-7DgX<9#^[X=?,N==Dd^,
;V0c1D,[N?cF5(@g^0&>aC^EHBYd0MM?UKXYbH9]F9J4M;g-94Vf=K/E+Z+/<7ZK
):8;2IETJE1&4B7WRAJ)6;R<V4FeBF.;8SP0NJa5S&3?.OHA76OZ:HT9[>O5DIZ(
X-#Q75^&_XR1DFTZ<-_D;FLS1eM+afa&NcbO\FL^IW+b<S1QE88S=+:aePW/g;dU
a8;eHX70Ng,579G377RYZB<HgNbW_Jg15>G)=&>(,[A0YH+QWSCA30IJL:\aY6LD
K\\HY+AJ4XIA0=EF[c_NZ@T;Tb)@1>_bL>MJQf_)g,-M3#]4M(+cS.W?FJ7Z<eMH
)I<1(,40gO)<,R5-0J>OUE6HgV2G<X3g\:aJ3?CVA/<I)G.OHY_E69#[2H8-Wf50
W5YF43PNR@NbX(U@2Kg58AP[1/eHK61[2;9PG^@c,c&H>2B-?RbV@;[?U[fP:J:c
.>fcaF[NN_db;1Hd_g0KJ+(&LO164?:M]5bHKH95=F1]=/\Nf1V\A4DbELfW8R/J
dAO\/E8^>=&=fTg+&DUA@DL4Ve>-WV50=V[D+7:33fELe6d;Z&(C#:618MZ\B-DY
&72:LF?PS,UG8ODFOf_/FOX1QfX-DT7S14a0)&P,?LdI);1d]O(@Z/6@1,Q\A0CO
e<Z2[_WPbaN+,KG^7(WfV]G.F.^&]+Cb/WF0JbHCU0XdR;[\Y+P&f\H#JLa=X_./
P0X.b4.P)1#.LF_O<RNTgaHD#<>;)9K,M,F^97+G#+#0]<bL\41XD.(2IC;<.:]A
+>MJ7Z?0O1^\?PU?KQZ36a)<S5ML+JFI<IeW^eU]R<NB[_>Y-KTHIQ/@QJW-)TJ2
=]DZYV):RXFILcH+@G=.M_>I>R6?+@UZC,EeDB&W/D.@Pb<D:a45Z2:U.S]E/NNC
]UWPgOWW0A\e:YLF)1HeZ<C2^+Y?KF=(BLae)eFGfYWWX<OW9=AIE:X499^.4d>#
(E^H(fY4WZ^SEU,dVUYF9)[d?=S2>[W7WG)3Y+eCacb,0-ZZ+U6U?3Cf\QKWg/VE
:cI4K6X3XZ\:,@M8XW_g<UW(T:LfFRG_@<FQDg@bR)bdODS/1.9U^+&FdH/]@W,V
PWZZHU;U5bN<MX3C25#5bE6+4I)P?e?NF#[Q3ZF#6?X+ZL0b3:V:E5C4-;RJPCU?
aO87XP8fePe8WP+E2VJR2NN:TQ;:/FD:>YX@=c/K\e8B@S:=JRZDN=[D1(CSY8Ag
P&3LCX0RB[U.Z:7U)(81(+7D#ee&;+Qf.H],2Ic/D_SVP:/ZS)-LC@SZ+FXI?V\d
IA_1fKZBKS>a,IM?+D845ONc>DR9#P+U^Q(CQ/::)5HA2D5c>NeNXNK9aV7?W/?>
?Dd@3?LD,c7d0#bXG\VFXB&U3>CYU+KPTB);bDg9+AWcKOJ:C\V02GFTB-QDVBaH
8c)17,6LWJ-[f66c[GK0H1gLge]&g2=2@>.K_bJeO#M0.FgFAdFL0<YPRY#]69d,
cZ9OY6#C9e4UC]g@(T8RRF9:\L3M.Y#\(dYcK?&cZI^ZZ\?0@H568P=]7>TNTCc3
(V#9;>LKC4eK\.<ZQVA)ee8H[IIaA-+ER@KA1E@MW(-SFS,<7E51HAJUdAB:+@E5
43&>HedLS#C.)/N8FS^_aR0D\OK(G7\0EXCM4S92^[;@dM9()G?8BN=8J;:1O7[5
LXJP)4Mbgb,D@2b+_TP2^J>9EA6#?G)MF0AE_gYSA=L26KSa[b\3V+_P?)U[O_c;
.FE/0Ud0N<]5L2bBbQG5ZbWV]-4Vg5=<dB&f0_Je3Y,6/b:9BB1^BDYC.P)/[S^B
COfeQN)7de\[;PU\](\SF6PE]YD].0>Z@I@XYG>]TOKd@<e:(P7(f#6^1:(f5Y=Y
^Z.G\Scc4S^39eC>O0I<_0#Bb=dV3;[@=]b2,Q=QJCL4[T2U2>Xe5TW-S8AQ45.Q
@&XYO177P;<T?BJD--8W4#=VZNc^e/GL>5\_JR.d7WeJYGZ7RUe?]W^7D)<g\#F?
=F8R^9DSJ02fPP7Y.Y3EM6P=8P0@>6ZNK9^6>J17)BQ(4]e^5:U12C[MfK^=UQGO
O+><FU#0bK;/&C2-#@ENOC-0/#&1XJ5HD6VS2S;WX=?E0>?BM/P,ZJJe)]441LXg
@(,3:_d:M)/HMKO5(-0B+_dHI)2>L5Z#L]b=2J7<(]LSA/4_f<PQE#R)I;H\Wa-4
W+^_Y0d2KCUa_709YR;<(V^XFTODR;bOG9C^^a@bMW;I9#dG&,dcbDHH]CL<aWa,
B?W=:DGb9<7M<,-K-Hg7IG.JaQCf/66=GDC4YD:_(Q\UV<<Dd67(),7#)MVF)WV8
Q<60P=.,H<,,?L/b4_ZY/3.1gQN-BGd=/[Z3JaD_BG7dc,c6(7JC-;f=[M13J):Q
^#6U2IC,&OA6[J?_+Fd1K;3(Na\_B.,a)9N6YRFAYMZFF69C:K8R#9#I3.F)IKC2
3I/57D3TZb75&Qfc@#(<:+@6K..K/5=GE)ca?/221>Q2(fdZ^PL1/V#Mcg[dT3b#
@e:/2e[F0YAZX:eU2WF=+bIV3[I&Uf?+Q[Q3^+TcE-VXBMS,Sc.Z9OTM&F;(<aDD
Y#OfH&]aXW=&,./U&N8fB3+QD\Y4O2cC=5CaC=RE(QQNcQDNS;ZTO1W02R[:G+C6
2]-L5W5#S\)7=3c>)GaKX<8X\Y02+gNMDeV6)RK5\0?U-C8:9WK4E\1b@D\MHc_B
PEVHfdDVN-M)6#66AX,-:+CQADR//+J@Q&ZeK[@TJ/bTgb>3^9^KA;NQCdQI?8J6
KA-K@Z[]Rf.C>?LH>,d.SO+8=62T_IJ@2M[LW@Bb2I^-C1_[Q46@Pec&;SPIa,_g
#f1a+:2SA-MdT#I04[B5bU^CH-5bc=:LYbfdWB(]<LKI]g=?41c09+a88+HRK6eD
=)L>Hae8S<Aac=ETS7C\SXOZ:?gb-/7fM_;@E-QS+Y@.5DB5bJ/#=5.JZC4/b[G7
=MHB<C#g7RJ]d-3/]A;#B2DR/f:K#7(0ZN7XYg9<8B<B0MY.JJE>^(_IUN]f,OcU
2/RUFQXa;8,Q=f#?W=?eNOHa;#QY&Gg;b^<SU&GUc89Y?/L69-37>=]:QLd,J[,D
:O[_gEY)dYS^f;DWQb0gOO5D;1b6,(U(A&]A2P]AXbc7Md>;NJG07;Af&Z_BP_D5
6GG>33>_XL/dCCa9^SW.FE7d:MI.0eHT[cP-J(X0+KQV>X8c<\=K3V9)a/SRP>U=
VSDZ;1W;(#-_OECRF-5fXPfW:-L18+&2Ze#EB?W&7X^[,62&1-g@N1cIJLU2^2EP
_D/13>]9]96SL=,K\P3C[KQW]c[&We;ZK4LJ8d\6>MgH+T3S8:[24>@:YLFa=32B
d<UOKWIR3L(O=&_<]+;1b_/8dZ]NA0&c9fB9f^JX4^?VV[_=YS2MIH/Y.4R>#Y2U
KLbRO5GbMV0<)73&OdLXOR1EOO5+M8RYWU2#)6^]-S4/,GDZ7fX-U_7cZJYc.M9?
\,C[#-ECA#c);<Z:]L<e,T[(II?2MD1M^]D6::>3>8[609EY:S\aWd#e]d=_a:E[
0(>+=E_]OUeO38[[.SG>H)?N83&PS\TTg3,9(1M(X3.),O][K]eE++Y-Rc/9ISca
[H(e:UeJB7cf_c1XKg8+.(a_@g63IU7JC;b80,IK@;gb,0U#M+X_[aMR?I0@_=41
SU+I==B_9.&[B4;]e1f>IL9/f-H5([=G52ag&d<<O-=0VTLANVa4R_:Q55M]&OBU
OWFSJLKU:Ha+e2Y7B>5+ZJCR(<KF4@^Q]a9FTa/N0D^@T<\EgH]5f9]9&ed7\XFa
:O>QJf[(L0A#F-=Z-PI-K1JZfCJ->4PIcc]01D(+4+9H2P#<Eb<Pa#/9E[&:TB]9
g?7]g53X^M]IX1AL#3cFeYbT;X:DQK#ZObW3?6U97J)3JcbA>4?YZUa>FCUF(7^0
90=#/-S?f3D]C;bX+3B)(D9@P@d/-;ITI5CdDG<<ZW<1dPK1=#Vb1B190I#(^7WS
5Q9&7AB84-=VLP\cVR)4XHEReO7]=9JJd,<Q_A@-KF0We,)?X68TfcOV@58U6I<a
^GS;>\=3&gZ(N0^A@/Q+N<#AWM0Q+B\&AV^-&T[NN.N<\g^@I521>&P,b4&TM]CP
HceI2<HTIEVP(A52e1Q^af=XBM20@0=>LD#0><75O,0Q2gI5V1]T]/T<Y:-?Z>;c
baF=3.GIKJ-M:YX6HfT03&=Xd\aW\aF6US:Xd4[Z?U7M4\4,9;ZG>)f:2d-HQT48
BQUK\0gFP\b\gFRU.8U,U^-O4QFJ7Z0\.ZBcMTJ(E18\,c?I^]DSe1f;6AVK;UOI
3CcbO7^?g2MA1C:T7@L59H9g8UfL72XXJc4M]f,,,)DY76IYC>4&3G,GVHZ&.eP,
BJ,][:2)KIaRZ30I^4^;RS68D(@S9Z#/BZ(^AIOTaM/eI^YI[Pc;Bd1(X,HVGEB?
:(9MBb7+KR:ZdCUINAbS.\>9S+&dZOGM:(&XH4,&@W@9<P=7;6.D]f7T6FH6C5<g
>dX)V)eX_W)T-HffOXQIJgK[A3R-be/?FZ:e>@\^-0@>)Tf\EN,.YADI2\=UT<88
(<F;+E>[S)U78X@S4@F_>YRedF\T,#7O^Bc?AC)QL9KdPYJXD3Xb9B_R:S&L/#_D
aYcdS7Bg5Eb6\TQLI6U,eU/1U]5B:,<?cJ>GNU^W65dNcR?HX.gdJ-K9>0DROF)V
,Yb^@N?##fXEDf&Of2T\U+KPEKOfY;J.X.^MBRg4Q_1&8O:VC8V09@IA7-5c-&F]
?W_c9@N7#?4eX-SPgC,HJ]A3KIJ>Bc]6a,agEC]M_\9RXUZC9JaLd?K1FIBa<eX/
V5A&B4cPRg+9/95A1Y0A\PS;WJMgK2W(8N2X+XMbd/:1SCEe50>UL:JW+)KV@gFQ
C=T/XAQ4bA=b6FA[0J#=aH@8T<^I2)]e88)c20NKfRD=AW.:-15^^4&1U0Q@A&U7
D4;]bBGGPfB>/S-_8<LQ-KWGIc_D(XSDHC^WIL6#L?>83e[]>a3>XMQHEW=T;&UL
SDAS=FXT]H[SO?8b+?LIN>25XE_Q38#S8NIa8RD.(K+DH9]J;E.?DQ2W(JP;RNZ#
#ZXN;QQb@Q^VXLBNS27L2J_<919ZQ9UN^>@?[gS#6ZdG>Ba7\8eLPD9I:/.A]KY1
4b?LCJ\acK=&b&fV+dL3>:NGaF05T&R]G-CXP[Rb5;=J;gU9/C&>P3NRWLAaLcD+
AK4T)b&b:_PeKPe4Z<N,OKbT.:Ed[[S.Tgg_4SHVG>Tg-e#QAaaRYB?3JSdUXLMF
D2@D:R?5_Og6fCe9)465CR&_c)S?&6#-PJVfQ:1_WN?YR+4CP(?=N5dV[]>DHeHF
\<3>-OBSP8(XGS-QZ--\6Ub\EE2C5e<,dKUUHZ/)0;HXFEO--Y\F,OUAE[KS(:A/
ed@1KRAK:\+gEK7+_+W7,SV8.Z@3>QV82&(KV3^]+H?bD\Ta\R374B#/;ZDY60F3
NP_cX].;Lg#R52I=XJ7</&JYBdUcIM0Y)e3]@T<<?O^MG@;67U(YNb3081ff/_)3
X,/2Ng1\JST(7.UV?:+3GMbWCRBUO9M2OK3HN(3-\bKT6GOFF..RBO2?378@;]af
eCR5GG&eND?^5=+.?1#CAZ:\acWec>K9-+0T[SIAUW8Y01_O+[ZD4TbY9>(/B;EP
;K4FFHP0B#b,=996D2_5/4_f&WLD8DgR>V[@Q(.M4P1>CD?Ta)6R#?420_H5DBTE
a7YA9QP0;]?=[;4MXIY/1SPf[S6d\I/]5Q/&X1^K2]P[K:;D_<,[RAW8U+a383JH
(RfU-)Rg9fBc3eBc?-9-Df&E85AJJ@gDBDeAO^ATFUcSFa//0#63_f)IgE:2eTBB
dC7\WgN@[>=/N2.f_F64>V#d@]FY<;WTO]ZLM1Y7#)f,(4?>)e0Zg]PTA;[9Ngb:
(f?>VK3Z7I&^E1d=VfWN3f3KFJ-J/(.=6Q0]^UWJY0)V4/520#a5PK)]UT&&;;HC
JU[f?d0RB8]NJDJQQddLRB<5(+SMV(#6,6;78a-#GVCgc?B1BIDcYP1QKS\V<?M=
c2T#5O&1IXP5^I4W21Uf)S].=IN(VCTGgNHN>Y\TAKc[#?[F_NQbA3EbfZL>He7F
)c[KAX4S[E2R]649UZGRZK\9Y#D_-VfBF[94-+2>cf^V8VPV]7/>2^QfPP(R(ZQA
26M^43@SK36.X+7_^f/aSKSf5?-PfR+P^b-ULO_&@f,Q:171g0)S[O(Yc(WAP4)C
Xab,-cD=2aS6FO6D8\7F6H.:;T[^Lf^&7]AN[LGK>1S-0X7ZT,9dTJE?7-&J36Q#
e]1NC2XgQbOe@W78G08Z-+-FYd0;[^4+3+.dT/Rc(KFKV?Ad=\/.I5\6;Cc=T_Ub
/J7/O,Aa1b(R9R[0H^]DeDU;33=W/U^Kge_=5/CKe_]+)8VEgU0(ZSC]<_Ec#S,&
),dN:O&5,;OLdAc[9+)+c+ZILa<[WZ+4UM(<cGZQW.L<^D9^?6BINeCPPEB,5/5^
dFWAcM2Fg3YbCA]R[If+TIEbL5P;T]J4f3;W(M,b3DbNWX,_\I=I+6AFMEO>g6J6
BE#4,:eLS\e4_:Y91.?7IG\[,XO65F8+1U1L<MDP7VIS4ZU\/.^B8R(S_LAC5K,]
[2+?G#8b-R>V1H^&e78?DE)^+<5FY;K+87.J.E6MA/G/\c-F9)1N3GRc+ZT^Q16&
TO:E+0=Ng3L/Z],2WVABHUY0546O/4NSC=_&/.ab>&Jg8(,./;FQB.0M?R,N@@UG
9Y64ZHcI(fB1<@VdX6VXX[G4:@R0Q^a]Id@aV>P+Z=\MQUA]B\(V9M,@R4d2HXAW
2:01TMY>,+cJ+..WQ_KY^[/bL[?dFO@C@8/6O</Yd>^S2b^@SgFMG2cCQW@/47(]
<g5-ce1/ML//eH3gQXAY9;KK-?c[TG.++4B\LZ\NE88ac#3S+E0dZV?I4_6Q5bA_
S/V2)+\\EAeGY93)GT96_D68BZ&T7N:J543?VA:XW1E^\/;C;bFc^.>X<JH383C]
<bXMCH37NOX_G^3b+0X_/g80/F4B2BWYJ;QN.TgJ6UP^T<:e+QUX2-\\&Z(E=9U0
g1[Tf.11>:@BZaDTCHXA?+9aI@-.W[Y^<8+DeKM91XEE</(GR#0S#)>g,<#.1[^&
GLR26+KMPY;?(3HC@8^JC+LNc#_FKULO\H751<C@MGN<<O_R4&E]VW+H(\G#B;]\
Qa22]IMM&[_?-(4,Gb-V9b8G=3J@4dLOTdc#@R.2_)(.-A-cX5]WZScH1KHTB);P
\bH?G[ZD6ZJ(T:E^@6SK0d+cQ]VFA^C>Af-R/JeC7^V);W]eNAZ;R(f:dD1F/S^#
8\QUeY>g?Tc0;cZY[(F4V526[9K#4JQBI.K60I:I_XQbY4.3CDWE;?-26Z2C>^ZH
F>^Z/eXS4X;PUeW6YFWWXEKG7.S43SMGd]@eaTLCP8C</R@DI-e^BFd80C60G3EU
LN5^<g&2?M2#6fE(ePV&_A)]4[5BS-c\JeB.+c.<7BQ6cM&J<]CP[,gC6)Q+SKaX
#&;1>1]35^0@aNH.VEg>89eJ@9_>??2H;(E8TL6-[P.C>d?H<3\&)dJWef2U\c#S
?/DB7Y<R0.a9U6eKc98.CcEPZ3GGc5gL9L6g;:.J#,HL/Ma@;#gVW&L953CO14A\
+)&-]01bL6eR?(XV\5NC)E+3<1KE@+g97_V[8:BWA_A4REN/a3)E\/7:a2A@Re_>
_O^P202eg<W\RgD=&(GE@[g7ScefN1DG+&U&S2HB(G31>PgX@A>6)bH0+FAR9@H0
C3RWd^^77H<UHS&S2>)/C+(Y<PMI>4B6E1Zd<@LW1\&:2D^^gEOPA3e3cOT&[YQ?
IAA3A#8I2;EBY,N]=>d]J7-_M3PUR&Sf?L[UTQ\+2cbX5YU(3&/VF3>d\4Q#MD06
)1b;.c1.D^/?PIDG\GA#(1,@U^2W#T^V)1P;dg_V?A)>+:9D2AFNf+aJ8V&,4+2B
ZF6dgT;5Y]KR/JHK?Xcf9M(ffDa]@7aT^gP\Y14G<^AX[@bKRU?)::MQH^TVa&SG
UUOe.SKW:)70V+HYF_>c[?4=<Bf59REOTF7bQSUKCWZI7cH701/J0PX:R1,DO[U3
b9LPGE61=K-TB&I_9N6Y+M^F-9;NL[1#g_CV]G,L?eOY@/4#cU^W3-J4^O9(#eR>
LLQE70NB_>496eLbAZ^\,A8cEfX\.SKT<<@K^1,M4=?0P,c8d-6X7,1^SMQI>KAI
WY<W>/T1#+aF0.W@51RSLOB0eEQX7C^2f0+&5<]/37GceVf(3><P>CVa#1ffG-e6
.cK@(P]bC?B67.Z>fS(5#7SDF0aFWZ[HK@XAMeNSU?;BVCdFA].e>?S:&6WP\?Hf
U>RA#]66Aa1=@X/.(>OR>?ONP1]V?ObH[+A(9#R4VKOS]&P;H+7fYO=PLT8IE\/e
aeV:5#_#e,YUb_LFaeZ3<HBOD>A;(4,;e(\2#8b7CSEYB<&&3=&54&VK)=BM\C#L
b)S<F3<RQB0WfA++0I1JZ89G\bZ.SZcMT#AJX<=_P4;DJ)W0XF_KJ0Z@/@3O6]YW
XbP^K\A=5A2L.G)6d1-?Y?9de;Z&7E54URbMOW]H#NC2(cLRL;f;#HRBKAf5FF3]
.A>3#D.U(==5HeaV&d;B=&^?dF(2N@GEFY@#R&9df&K33HR_cLZI.[C&#b2fV.6f
WA@a>XJAT,3/;S@]b(_YKCX^cd]PcCeB?VKX6>7PP-(1LFB]_T>/U?O,,D(Y;AGD
<TH)=cE8URZ1TGW7S[8Nc;>Y/QN44#Rc2A8R9QEQ-IJOX7EHV0+JQ7Ud##e23CA)
1aK@.4^^T#c[06ZH@7dF3HSB,#2LST#bb6=IJ2]?W6,J\Q/9&aecbY&EY@YH6CG_
IH-BJL.g7)-HRA2WCGT(Y4O^)cFC@J\gT/=dQK:TC:;2bXU;cL8H[6VX799dMP>0
7(^>UJ<a@-f&bHRU-1N@1aFY#C(#_/L,ELM:Oc_3973)IF4aY.NWDd&M5EA.E6SG
F)[^C^ZS/Y1#LcLMN2AW7<OOIO8#+PYRV8K]eWce;R-+SI66YDDaSWgeKD#^3(bK
FXOFSSPfZ200#I/QIUS^QT-G\3C6[cNAJ=f^eP\J]5PX;XQdKBQ)#TbP1&I8^7Pa
C97_R?602<<2gUD#VKe#\KZAU\X9QHCD-)M+\XI)Mc<:;VM4L(g)R_=<RGZ&(-?]
?6HCc6;#R/+a3&N6Mf/[P.0=(TLXH\CLC\9-N0WL=LYBVEP^]9AGP.J2YN<=M\FG
WfD60DSfRUeFg.LZ\:\S;]GM7Y=9e2@DKNP5N<[,/eSF;6OG=O_[.P8d[949VASU
cD7C89>6?/2f[,]3b>L4GA[MC-KcBe+K7(K/G4LD9@#A/(+/&A.cN(UbZ-R1BYbZ
c5g1_\K0W\SOMg7^<1)-O5-NO:?YT2HB1=aNJfa9RObO(@G&8+TRV:#(U8>GA_b#
@[a49N+>RJY;fbfM^1Md^.K);=#2YFVfcLJ:.46Y^<V&1T2YX_TdN(S-3D]:/..b
^J7]6VEZOABNO&LK-GH7<KFP6[>9W=0N]_2#&NE[2-B./:HL6P7,@D4[\V1HB#4/
[aPY2?BfX:RSNA9(L;Bg\b.d4AX=;OI3?\cV#ZNV6)HFS+-VWJWf2K[FK03H\U^V
=T7/QB7ZG&.2F2aOM>N&)AObMW570+PUMdJN[I;b2MBA;M.9=+342#J[UY:E\:+F
AdHFMTM_,4Y__#)_Xg<L<@9F#,N+aGK&b,QPgTFU;bg./Z^Df/<(fUeOG2O&YC@\
-1OA5@d;gVKYcI8-]&H9IQ?gee99/=FVgA<P\#)AI<@QMWcYA:8Dac4H8L<;)0ZD
TfO0QEX_JG,a5=a-bId-a5O-(2;?3ETOEcX?4VX6HW)<TDc06_NX^XX]FP/+5e&)
G)bB?#59g_36gKUB2e:/.TA2CI]+d<6gQ6agE^T&JA:6G#6+7<6N\G&))[(6T?Lc
(/M=]a_CXRV99-R=?2RE<\_EW/4W=P3:C-X>d5^?I2PZ5N+,C?=U+=C7D=+_81U+
Xce/>]ga&KQV+:BJB:=>JKI[SP01\L,H/?H+4dS+HPHP5[#VGg5/W+V>&U8\C(ce
465WQ\9=K).7Q,.GJZNX265-QK:_0A)ccPg[fH4bb.R,+JQ;>5a+Q/I-Uc,f?X6A
6_AS8#1N6#fADe@KB>HN.;3@/B]W#4CW89(7CV?+X[3(V=d@XYL;Sd_ZX)D#_=>\
Z7gYZ=02E@B4Y/b)G\:.]2^IJ7B[&_<?6E](7UYWT@,-a^QL)RDJUTY;9Z1(6;>I
>b9+bf?OQNKGMILM#KdIYC?@M32(YW8O(WCf+X_>N.EV&[\Z]YDA/])>=-?c&d^9
6+9-Z=D6UE[60W?E\3/F4X@CQ-U2<):e]+UTO59@_5Kfd(D<M^GUT=KNVR79-?[I
V&-U([;^/,g,c-Q7f?JXL)S8cE);]L/+g+bOGCT4_;(0;A+P,@5F>9@Ka3YDDeDX
Y[(&5]9-@X-HZPU,8dRe::DPU5YfgL7fW3ZWE1N92#ZI,,X_XLX[V6Ob5&PgKFJ:
]U<BC2CC&&-ZT-I0\eIf-1/ba75^8A840==5JV8UG[HB4C@T_Q3D<5F,:__V?ZW:
5.:7,=/869DHe6+E)=W,Y)PJ;S3KD&/N2/8?afV<BDS_S:#aJYa&^Z5JHbPJ1U)X
S3),cW)LPd#.P-(RdE51W4TJ7QYO?HEA4Gf6g69(5Rd[dcKAf+RYBX0T:Y+=B@7N
2[ICE;>\e71Sb+Qc=[KcI.ACNMDSNQ+&g5Z2<H;-g_R1;HcZ4PG@0Yg8Ha_bEJa.
JbGK\93P[A;NNV[eZ[1CW.gcC\\\.ZCSJ2:I\XW_QR_2.ONf9;BGb76fZ)DgO]G,
-S8^RIb6FQbRg5Pd)Qa>13M_B2c+7?@.)9e;6JI6LK&^TC8I?LM6Ib^9f1.TXaO@
9JEJ-EA_CR<N8MS[QRY@\1/2d:+3#G_<g3XRbG,bL<]79RCRHM#.\4&IT;,5Q<AK
]6)IPX]/_(1cQ4I],;MeGWNS\\:NB=+7Qc@]ba4KN(F\PY@5N)&Z[C[fe6Q@,#+]
fFMXK:?3HcN9<eC5-8QMX;1(+K<;P\_/1;0\)_DAE<T&EL:X/dB4PYL+e\(#YW&^
:2LO12E@FZ)_-1f8(1H0,b0AMNGMQLaU0TQ(FF04gKW]GM8+a<80fX?+0/HSS^d?
C2;2+_ab\GI+7&Z<0=g?PEXGZ9<E]6[^I?L8[/a/J\)FUET_3JZ-)G<-\N\L2P6H
N[0:>N3(F=BHA_NMW=&_?C,X(F(Fc\e08Ve2R#JLZA>=Yd,FbDc)XB]eAQG7^T+g
AWW/SU6C.d,0B[UEFNQKSf->XN7Dg4]9L/S1#8L#7+)XfTEJbB#@9D[9]I#1PI,7
S)D0Hd/;J5^BT/<\W9ADH6O?gU7Y8I02[O4TZE13\6O,+/._DdeWEN^L;\a;EZ7F
KQ8QJFG1d@Hf(4[1T9S:>-#cWD)GM/=H4f/QI43-WVT<#cZ7BTgD/69(SC&7\f;&
=.--FA-T.2f1QPMQYQWXAFLCA/+^.M:6[;PM(dV]ROFH2GUG@QK[c2I^JTcS2ZNL
)^cL.B04ZL,C,M4fJ_?_37=/;cCX+_KPM4G_94?/@I80SJfA1M7KZRN.?[D>Ja5#
_0I.a^JWK:?N>-C9>JY,O9WeG3gG/a<a41:B\P^_2aO<VXQQGW3=)TV?YUV[4Vf2
C?f,[>c;+7;IWNVeA,+:;]dG?0(3)+2a>ZU\Q[_6/0fM##4._0Z+R7V?eB)=(8[=
3TQ#>M\([<e45E)d;(KS-R0AKb6bX7e_E.51NLXeHe)>48\;_R8R_8>-a_H4ATD#
CN^-4@<g>)LY9588DgAb/RB+/E51/4+3I=S>N#UdEE\S(H_=/)VS/R-J.,>^[W/N
^N.O-Oc[ONM3??f8C^JG5LI6KT^KLADDY3)U<P?]e/)3N0&N2V(^HA61cV?U_(.I
6V3AbWF(\C_VHTe1LYVSA;H96/J&7>]\M[d_[_gI5g2<#,/&=5BPBJg.PAB2K9d1
935X9IF+GF/J6Q8S(,5Y<@O]E-?(ECP@=:f&.SN95MY&E>[?e^P(U08J:@7YI3M4
&?H>)cfB#A8L18]7=&M6fMeD)c7fKF+7Y<:9Zc9I=0Je=+#Q+.@e:@]GdR5Ha5^4
V(1AHc0aCSH2Y@PR[_6b]MaGcBH88e3cgX&EM_P\X#[P^UHNGQ;A[<[REeV(]@#4
4^&gJ0F]NQFaB<1X6VAcH=&cFW.0S7--50ga&6(VF+POZQNU-aVC&>CaZ+X.G5\(
;Y&ZEBI]KCgUfM?c+_2/f_9JVD6:1d]gZ/KLC(-bM+aGNW(Q[77ITT]FJN(QEB:U
S<CRH6c&.)NH)eP[AHaT,:_+fMbQ#aDcPH0NWVYN#I[><2A/Y2e=A8gO[;NDIbE0
H]VSM:c01?A3cS;NH/E0a.3QOKVaL_8?W68/NZ:-HAHCDLO?cNNR9ceB18\fNADU
;-La/\TJ.E=L:L,-ZK,>??7?_01Q7baLPZL9W8,aGD9F^deb#GJZT3>=8/ADXS71
>@[(E;Qd1-^\2,6J#IK80HGfQ0>\4&8YT01(MT6QLb5ec3Y<U2.d<=5PL0gQOWa@
BaMdR0C^Y/:W;F1C7URe]bX;.5=_Q)/Z9BdV+,J\M2MBB\SQ\@A)0<1^-VM7@WHP
W&F[3M2>4C\[4]e56L4PA1+6VX\H3P=4a6TV,GR6X9KG=&XANJHH;B?fK[@X1QR:
>2\-L>DIHA_ZYIT8E36/43^H=I]LZT#^^X]@<Ocd<P9dcLE21Y8GfHL[_P-Vf5(C
RdTS@^@ZT?B<_(8REf(7LT<8I6/Q(71:ACZ/ScXS2KfC2OXIU&ACN&FOQ1>1(6,0
K\SM[ge3G2QZUF#U3c>FX[H]?P,N-)OIVK^YVQ/H+QIG57[ULe:WbK,g8+D4H.C8
eMUZ[e=TTX#F]-6MK7@ca<D4DL)@@-8[DNBXB?cRT?eFf?I5PZD6PT>gbYWVO,(/
>6<^27)+;.TKdTTbEX<6D-Gf(f9Y)G):M[>+<>;__O^?2-^aB]-Kf,bLG39X>H9O
#R_D;1/72H02gHa&eSH(4T-.g/A2#,ZT3SRf^/ZM0@3PeAda\,Ee_\YTGU@(C3gV
7J=+2/[,=8a1P94-/>;HAA0]B5TFHODC2?QNG0+3K/:+FeDcea2gQ6[#>4,+\Y11
gfI)JR7PXC#,K0O6;UZ;EN/JfTRA-CS)PdYF7F.5<)^S<L&^gPQa8(?Jca^b._;A
0ab4SW9;AfPLA=\2))Q<^dCKb#EB[2GFSCW]9^R>=QWg?9;U5Z6(TCO@W^OLDN-^
FDQ8,ETfD\C-@)g<DC+IP=CCXa44MaP@U\?9X8DSf1d=CXS_=:eCc7Z18GCND&PK
93X0QL8=)>Rg84;,#4P#H;C@gDS/W];Q-.SB\51>^HQeVLc75SJ-5cMe;N4]()YM
9((?613N(3J:;>,bg1E7M=4P>^1MC)^:)DZ\7eJDVP2R8Af.Fc7=MZ2OU]\7:-]e
Q(8WEMVSX21M?E:BKXAF)X@NT)YNL+7HINL8;OP7VIXXM)N0e1Z_3<5QK<[D.Z,4
YT/<aW?P3Z>9@Wa):2TKddF@2UHF+P>AMW[cNc)90,\NC8Y@=<CU;+[3QA0Tcg^E
W;7aCJW78P]2E\.XE).W.eA?RJKXB6B3:@c\AQ&V]H/H/cHS8gM26-ffNcg@?+8G
6f#9MP&C6/fg,J(b]aNgH7(RKfe,:#f^<aJ-X?\9D<FQ?<gKF8cD>+.b8:Jd/0F[
YQcaNYeF^.d\=Z]E52JbHL@HHc#0.771#5HJB>b8Wa9FOMVGF@4+JY5>e4E+eD5:
29M;Y(TF:).84B/.^g9C?<<SSP-]0(M#12G,+HCDc/0ea-Z4a\K3++[Yb)RGWF9O
e2[a2+8f7aYX\M#+><,U\?E)XK.KB>77^ZNX8,28/fK8CER29:AG2_;U+PJI6<S:
@O-UZZaM(W4GdNN\;>[;/BA:VfP4L>XV.a]#.e2ZPD:&-INeE+8_Wb9RCIN[&>]L
>&]f.-(g,1O855K#VMP;]8c12e?G+&]Y1_)(])1LbA-Lf,a81/S\)6;dTSU_Xf6.
U1IOXfHGOfbNKaeO6a5KRFHRJ;MP@I1YD\/U:<+dH?CDG-JXQ9g,62+:fL3QIB.(
WX<M5[Z93SP@d)cC[@,g?T/08d+acdRG&>M&,b@0[F(#eA9AaIB4F?<;KVgC\^-P
b_CQK6I/P@SD@FJ6+O]]?,/^6d.SEFVDU.IW0a];^]<Z^1TQgI2;W:6DDGW8WI.f
@2#IY3f(cWJS(PWNI3fPJAKcJf2I#9bX.8(K,9Oe(OZ>;MOCY0c=.UIMNf^R+)5O
[7Hba?E4/UPTVHb]KDOH-^N,99__gg)848>SHebF;2<V8,7WBP&)1HMGW:6:?8OU
/957VK<\9X0e2]I&4.5AJ_acL/@&&HU<8T)XM]2c3H\[?N,X,;V?4I2UMV=50WS:
8C\7(+6S=ZfK1TJ@O3ACC,9Q&3\F1dUVX-e.@=D2e1Y55Gf;:g/ceS<gK#D3_2Nf
:Ka(ICea9[[Y5[]fg6F&T<EeI2^IRBQ;F]+@A+7MD/.Q+)]Qe-->/5GZg(=>&Z-R
/]?d>E:XfF,HIc1+?(N.+1,>P&\+:c.JEfF[V5/eS6<D;:7?2@,_X<784e+<SLY9
&Y[0X<,.I-Z@6N\ff0)>2,MP>J_f1XB7?F__4IcKbRE,0<K(JF]HD==T)Eb&c(>=
BEM-XY\>8)DWIR:Ke7dM^_:BU8E0OM2@.X8Kc>]/e^/]aTWV(D:.JXG7@P-7C]CM
T+e9]7UW@UHD/TSN\J=gF(IBgXLG,O5M)aFDJO_J^ZOIa\<KgY&TA0&\:ZfKFX>U
e=VHe2;S[]Y8gdE/QM-+0)7H9-U,-e<FT26^@.S,?Z=)1cO?R<WTJ9ePOW-Ic[<2
=54eZ74[aH8-IEF:0+KRV0)(9R+S>Na8;Z]GH_b:.Z?+#eDNAZ9N9NLI<TQW(QN2
cOXN2W1=LId58??eC#DDFDf&>.a:]<LN8CF4D>(II\HBWVAV5+LF@a_f9Eg9@b(H
QY0E]2cP7Ec)_D\WVQf<W@[=]+0:>J^(.5=6O/7NKQ4G<Dfae&]/O>UY9TKdL=<7
9.9ZbW8\C8C:c4S&E\Y3AU:0&U0BZO&F^O?deJHd84:A;0+b-7NT@9.J2Z9MPY\\
=/4&eKX(5ZNLAFT.D@=\A3I[\QSG,JDXE^W?^P3]XdVHGf,\?7;:J,:EK<7(U>^W
:K[=-4_9G>&(./>1NRR)46:T?22IWO,1aJW+[Q^PagGd/U,CTYLWO7PGD0-(VFUA
Kd7gKP@/BL1CSfC_;b:1A)\Q&NFWTW)5KOe^adOQ-F4N68<VT<B]:<7-KT[NM;+J
c#6eb\O><F<AVE_]-5Q.DSSLgX-,9I1b7X50aAIQR9IV-1,242)7Z.([QFgc73]@
Sb[D@?IF&fM+37d-:/Y4>DARLMY;gT1Sfe9&a<OP[^deD07-dRQf<2+6W0&4?P&<
ES0D\IJ?.CgSXb@/EX1d(TWQZ5J.I3eWDL.d3I#40I?^:)^#9=BM5OKDg)Q</:?b
Q1BYQ\92XNL9.M9+Q9@2@e@X,.8]COcXZFE(DYS-O0H6A3g>:/b,XTfH4LKDRMdQ
[Q-H@-+5UWZ0fdU8QNLNf97X+cKe]>P7SfPU\3BE.Y:3eRPQEA,V^@N<La,OZ0d(
BUZF=LE1\^ed&KH]b:\MDH9DBgZ7c^dOf8_E)6BWDSLa5EB<-)+WIGTeScP6;/M:
2I39+A=-<WW,[9_\HUc(^?HU#)-##7VQ<>)6VY.Ha\H;[^0??3XY+;]2F4L\BVG_
99H9-gVG4/a<aXD+Q&U1<RP:W+8U:Z#NRR>=?A^.F;;^a8ELC;\CO-d1HXT#\f3Q
d;dIY:bDPL(DBKeZ5&26H&HX7-d2>Ba0GYP8:_JW]J)Y3cW3Y,6a.@4=3GgPCK\<
L]P,44.P0G\)+X#3@1<57c@SWOR8OM.>.W(3KMcDg&(R&CGG,(:N6RK:4d;]7TZ<
+SbOUfTOI[La)X^aZJ3NZ.AMR5T.;R)1PXBYQ4MRDBK/ede:fgVY;;3W0SG[G]db
;<WfIU)D-P;O#E_.?<[:R)<W6,,^-LOLH<6XR:@3TU#I:S4.I;I)FDbDcSB6]NS2
gFSSVVd51@JQAPeXJ>>Ue.gKA>Ba8_V_?2e9ATI7^-Q;5<@Y43X3,G(4g45JH2I2
d4Ke^,F@Q,:(<>TN-2gB(cYSPQMeMIgAWcY/AEED:K3VQ)NH;6]@B7H7X&5&<MH2
5dOVeX&1;?@bDFD#+&a]8]1POEXC,,9e0C]=&+J()c^;/,H3_HaB=25L5L?R#eGO
1LTAPG;/5N+:9?ZV(#5OU1DJ2@Ga\@:RQ2XPg,EF@_/QTJ18O-OKX]-SJZdEd#=-
Z;KLWP<[P0H+Q&g.FU/6-J6]94a?[gYOE>E4J?3d4gg45HZO,-c<+6/1/QM5SS_e
/P=E1,3;-?@ZV;HB6LWD1;+N0>WE17&9cN5)U_CL4=<O@bX7=OLLHSV9U>GNK0gR
;V/9Z9.2f:L827E_HVEQDVBT5.;FO)4\8?<A#(_E)SDQI0F)U<Tf2a&gSYc7&Z0c
dEcM]>#GUba&QVV6ZOCJLFV:\N?YAdK^(R\AgE+CKI+^CI6\>@;8Ra5PfC7C-(d#
UR&Rf5a1gW<^2:2J.#G#^L@15#W0>N=eL-[PT/9HLdCJ&1c7?4,N4/PS/]-<M#dD
>f][7a8>]Ib9=+:6G@:D3V/[SMS]B[GDC6aK_?cL]@31]Ab[0M9XH@-QbPI)ZJeH
KE^L>433?16R-Q8R^IVK8^NQ.O_/U1cJB0IGfb[&B5FWFM/A^)ZQDVEUL,N@a0^W
K^g[\A/GA\:-G-cFL=89De[1]?LKK.M:6#6;M(O,RZZeY6aaYdF04<Z74,>8ce/b
@EZL2F/b@><S-94T4\)R\SFRI@\=>MQ\eB;=T/G-U^BQHG[30:>EWb9>IR&46.>P
:;;HJ^_2JOPN5HT5WFaLJWZ#_0,A:)?AMT#KO4HFLaKIMC#S0V-9Sb>VW8WG)G?.
K>B5KY0;0_,0;.1J=?=&?>RgN[_O_LJ6<:(d-[K;8J/3SR9U;Kc1I[B:_f4\DSgR
Ic#c3Ng4).BV&:@7Mc]PT9ST:N./3M+U32O_DSU[][WYdbgLH9P)5&D[K;BN:EJ/
&R(<DNNcZf\58Ubc+WKO]I_DN(G[CKX.R]M_/:@JDMR::AZfb6_N\SB),&)#V\[d
62:UB>2d0]VU^b&O@CJGXc&;@TFY1C4&;PXHWPIg]YJ.(5,EZd8A6CQ)cDC8FCC5
DXN)9Z&cF9QW#BAM&#XLcV1[YCX4GbbL>PEfK7E3L3?WP54_+#]FC7?Y;D(Q4cSC
OadbJ,=@Q<WP.gEV6>d_]J;.DF<>3cG]/9>(&(63-LESJ.9ND&@4(--7a#KO2I)1
,;_K3TE+R4U+b>c)3N&?CP_GWQQ6ZO\OXg2?4dXZd\@fS\g^#Fc(@2;G_^D=.;)9
JDQLX+VeW[C<bOHN5Z_87CFDZYe3<=H\1(cFUA&O\331fT)D//HNGRc\=VX+6-Z9
47EOEE?EB=PKW&Q+[G+T)_HKHAAc8f3=[,]I>VDY.,TfS@S50\bE.G=.\R\2\86f
,a6/238JbHQ7HgQ3e=/EGVgN<.,12Y&BXQSY@7,DFAZ1NY\d/,WA>MC]BP>M^W41
?9(C;7R^f-D]N/^=M[[13E.#Pe=1.(CL0W^YT(-U:=2>#>\N@3(c),e=fc2U/.1=
-^@c_;2]JT;QgWXYE(1SE@dP->77ZV\YN6cVa:E_XGLd9b;YSa0,/)_=/HgYN7DP
aO6)d._74:,&Z1(94O?1dHa[3cL51GL=ZYJYU4EL/OJW]=_ANeg^I12YaX9XU+=>
\@;UG&W#MFZC@7=T_[dTWY:@<<);?&F,PZW/T0R6Pe._&GLAPS-;1@cAM8Lfc.<,
+&IMGHWT6VBH/VHPXfS.>R[?V38=?b_M.3(_&U77e,;7+_3;Q1\SePM+1d8TL=95
SY.<U)YD0T#M<<>@<0#^1;2aKDV^_8>ED#f[;,^De.VfY)/D#AN\W>L+5@.Z6OP:
_M8J9RU0H?50WW<CO6+fBUA3(;0^;N;/S^4C.FId7gcP^-a]9g#b=?bZ\?EX@1>K
ANU)@5?EY4(8feOTL.8<KW9g@>,Cd7M]0\2:MWYb2_XX[6W/O#IcWDE04;0P@#K&
IfC85+KE//+Ud&eS230[cN//b(5RK-Z4=dG)D36YAR+fD[1G39JF(64TPC5H>4^@
^(e,/2V[g.+ab?8<9[TNWX#70KJTaKbTdC9.OX;L3+\^6B)?T\)<Y)\&5e.Vd;bE
E3X3,6<<?J;\.8S^=dH<ELE06[XTE/]OB0VQ9QP31K.@V,ZG/9IE@@7>)96\M/(^
UODNVaV?e\JJDg5>D<:0P?M^JLB;;N.(P^#DYMS2=EP_/L6f=;1U7gQDd-@.M;=-
[ZH#YIcEcM4c-W?6A[:(?d?/P1&Mee@@VX]dea+U)WaT&3F[V@I#P7(9H0QCdd15
GI_\06@ea5B,+XX]]F:_RCK4^QRT8F3^QWBGeNMBg<VaEW4XRHa>E,I=N?9H>KQ0
;gP:b.;HT5::,Jd1OQU0]=R)@Uf:H;Y(J<-38E(A?C_-9T8@Y4TU-G>-?_;TT@E+
Bg571/Y2.KQe^W<M88K59P49-]&#PY.S6#I_HWfEGXYOX,X/eeNeU7_[f#;R)V/=
M4KWO\7YMc,(:ZT4;@6_a#(8aOT^2,7[RcQ]ebO>E:X?cR^C]^X7@?-dGF58f[L-
c6ZI;,N:V<dX\13:U^[H49_D^I.]AJe...\+R_6U<3[K;-,1ET_&0;U\ET\9&YNA
a5EE]=c+VN_f&e2<G\607QN)I8eU<5;(QHfG56AZXW?UYQ#eDN>T><EBcI\DeWEY
KAGdP/GS)F9GE6)T<S8eD1Jb;1M59QYW40CcA\6BVM^=XV8-&-)RO4H5dYb>V5VV
:PN,LO<OL96ZY<N0Z/2W,7bE&C#04FSDBQJ^8ZHce?<K=QB[&&8Y&.&#O2,N\&KB
U\)SA4N\MA8S_-.)&PESK+7T7FB08>fLd_FXa4Rd3fBW0X]3CW;S0_WADcS4(df&
JN0T2TRRIZJDZ:gM57T.?G1PU2L<G]UO(\X^=]2:SLdd;+5LIY^M)]F@YG1=3G&<
Uc>YYa>d[@H.a7##fgQV48WKRAY5gR-.#cPb>@Z127(U/>b,,O?S?6H?c]^J^N.W
VM]21Qa?.3Q(3;VE>b8CA/TfCLL<@9&BOU/cV/bbbHQS#HO<EX]T1>N?3[=,DH<=
.EHC7:>Z?F&gQZ#;]gTDAU;.:R[J=NH[\,+[Wad8D+]&96(e9+O+O;<OM)K2Q?&M
IDP_SD]g?&BV+E^Gc/1\3TW,7-RgGY6F+>WQ-#+F/PXIg?D^J6#8[gTUD6L-HgF@
cbHS,K70#8bWN1:SF[A9M3F1V=XK^>#BDY_/XE.3/XWJ-a]H&g#7<,741B<g:I[d
KV&F3/T6/dQ)<7:9<,M:MK]13eQ1>SMFAX=(^I>^\>3A85[D>BHNE3ENX@_W=T)X
0Q3_;E)-\]>/YPP,7c?6UMe.b=ECG&K@TO1,Dg7+F6>XW?A6W27>eOK\HEA2LZW_
I.+bU.U]g2Y4[KO\Me(-/9?.]Yg:/:3/4;_#c899K_2:3f4VQG5ZPCUK_Vd4?V)X
2IfE@7#?>#2_)533>B82I2CgZH3;2T5)+PS@?f0JSeT;<)W/A\Oa:(YCMHO0HA5f
,6g920X19f/X[FNDO4A/GLJ3@7066@fcc6L@:1<BLW?AQR)+UbY59b[VPZDCPbY2
V[1058^J?=&<Pf76T=EX<fE8G4[&9VWT6V&aAYH_^Y^2V,__-E[DE;[e&B3/V7I[
-_=<7Q5cQZ0+53fUCQ&B\T33D8KK2X2PE<D>#CF_B,8/S(X[_6[P7(]RUf55\)Xb
IOK/0JIR&QTa4@<Afb92PGF:G\8#)G/)95Qc6d:GX).XZQf6B0B)-@V9@YY\6T[b
:2(d[<Q18(_DS@2XUQgL.#>?#8F;XH8)<>HVKf9@8BZ>@_Z\)OgIL+?gGX:5YMR&
\CQCICb[&b(.98LA<>I:SWP(Z932C^PYQFgc_e(Og]_T-D^\O_5Dc6_9BNVcL)-K
=]WSYC&2-7>bQ0d&S3J96IS80e(K:A7KVNDINYM_+19P2BD&fYcZ^=OX5@gZ@/85
@QPCg15?bV5cJ^ga#cB7&UdJ/fW^9e<B(35DBQ,0W2E\8+NLDeQ2)/\b1@13Y3Ea
W7F@B>+-[5dSS(9XEYX2;NA8Q&=-TCU<=R3(1,[;H\UT=58E\DN)1X,dK>ZMDV:J
f_Y&7+<R3:)]/gOgcg^X<AXLZWVJfIf.2.+]546T;LB@7RF]I0+,2#;0NN<7T^@B
E6;78_#B1CE?,#_YGc8\:4D15)XLY6:&&Ue18<Wa#C)XbeHR7QXGRd#2F4[ZQe&F
MA)fR>[,LG]ZB^AY-)\B5),@#KaFZB500dL6PF^AG(/D>PI7WR69b9[#GU^b6U89
=9Td_K>75c5)L95XAWI(QHRf&57V?<][=9RT,3X6[MS1JCbTK8<R7dKb<J-RMeVb
BbQ-FT8&GDO;@&Z;LY]NTSV-)-=AagQ\@0TXE^,Y&Ue2?R\H0^N&.aPA242[O+0@
;K7RJfCI;NcWDbOY>S-DP^0YIceWN\M^T9PK5)E.18^2V)d6B&]c-P\[(G^;UE+F
/V#?e=E(6<(QM@2MNU^4/L5E/#K<9[2?J(2GZ<R_bU]DJP)@bd=P;]bP_9(CG9eF
SUXH3CDgFM?VU6EN>T(;KC)7H0Qe3.bD,BV<-PS_\B?QGRaGIf3_4C3R07K,X)1.
8IH-?6BSW8c]H-&-[Q@)M0[XNP(1&K;.Ya>UMQ]\NQOC]9HK9MO83M_cNRWCPLX+
<0Bf9T?T4c>4D@aCSTN5CZV(]RYO,H8;K0\[>M>]aL,F\<LK\TS5;;>aN-Va&2C&
d=A\6?<Z;^RO_<9SQJA.,/N6J0;I6DbaN\&T/_:?WO[B<EO=DAb@^ARW@7908@bO
?+H8]NAM<U6d)X>U,.PXgE#b4P=V#&ACSB/]JWW4^A\\?B4^C(=8I6A,&A8)6)&6
(Jc\#4JDVg5W)Z/#&dQ(I4L>24T)SeVgUe4P&GA>e&B_3?D&]B[W0>K_6^?f6N,Q
JOSe-Ig)/I^=EDTV@Y5=QV-]SF710V.OFHUQaPFfb1GcST.Y\_OdCb/31f+<XSaK
eT[[QFbS]:eT6OIY-CQ5U&.eOPgQQRYZD=dKHT6S6?d_#3,2[M<]X:b.SJa:,Pf/
Be=#Ia\IVAV8](f78?@V47DUG>CYb#3dR.)0G04]X56,.&Q6\A#++=2X\g7bOR_K
Ae];U0TQ-Xe<bEX[8Gab?-.(a0aAcI?8g9WB6@&_^N/MAf(N1c[KK6E+6#9ae;2:
MO^dL[J^gM9,-7J2T3,BX1GC?@bb=SNK_4IQ77b=E:2f6A+fX^CeD2QZGUCY)#Ie
2f](<&M;,VFc@>S#65b,<MJ\d>@@#gf@fg01[2QO1O3X+S-PRTY+V9#ZVQUY9PNf
W9@S8=56]^UfbRP0+PA_K]U>6U8BA@Z:CUE#:eAV62JALdf@4AU>AO;W4+BeI0^<
2&THQ=1L11DM9U#KK-,gSQN);c@27G?<I8YYOg..+X/S0W::ELa?.]I/.(O:<5]a
RH0+ZFF]e12acOBVZ+aX?[<-G?F)T2JYBD^?TJCQdSCD@a+c>SV2F:g?&,\W8T_O
W/LG-TV[b19.?=8,d/]O@^=Q-6-O4:@2)39F_D]Y3Z9T,2?O@ZIQD_2^ZF27OC.C
;4LRM5FgQdA-/H+K^MeR4\M-P[&F<GdE8L(2/^NdHTZ3RI-/\d(X4,eU.\MF1d,M
NM=W:R?RKWS70Qf>d0C?+R_g=4?D:(M(I1N^aPD_)\P^+O4ZT[UHBPIT&F^aX[@2
Q1dSCH<K;\Y@NgB]aG9KY-bVB2.<da#<@TABNT6PdUR39^dE(8A<;KfA3]U@@4^7
88X70g\U0K4(H6OQIa\J3T=,TU8]ZLU4[:bYY9QC\2S6\a]24gEO#)J^RZJBARSZ
<d1BfA2RTTZ4)8Y=UWB7/;IPSH&:4#>[Q+Z9b:59_KE.\Ig@Gd-BD[2W._8K^<FO
S:UNc\HIU6b&(H>296-4:ZGX^EcF-22A68N3.F2N]1C@.B2+;50TG@^C,6&,G9#S
3H2XH@5B>XFfN)?-Pb4G@#LH(>BDS)Og@Y,Zg;7=>4Z^VI=aNEC=:;3C<[&MY8A[
&S;MC_PY)f#Q,A-_\U.3O1Ne#TfO6QRM4.a7@ad#_cV[:/N0gJ;B[06;&eWGE6&]
cf=B/Jcb?ZLAa9gHfO(/-FfCWGS:9.;E1S]+K9L@XVM(@&YAYWO(a@ZMHaVV]3YE
):HA9+bV1IgD]-Ee/8/KPMZ<KcN=QO\,LO+@Q/)H?X6/@?Z/3CXGbf?JE<L@#119
I;;:<X)3V^==;]58cNXD]P0Q7?,XSUW=0D5b5V+TC==4C6N9I>>MC4=bV=a+2)PP
-A_]T)JdJK;P8PA(6I)FB>g_@H](Mf3I(#/;Tgd8WLX0:E60bEUQP650Kc#L;OO)
LdLNCW5J4HWWC6<=J:Sf&34^:]>M(_4AE,L(RSAaDV(0I2)CgP3Q:(POV7+b22ZA
BEB&I.d^G9H<HSYUXN>,D;6T_FfAD&17CWRIO5LED\V<5Ya5]>(=\U.COZ[E^,Mb
6+>XRP2e<)[;<#D^OcZN9NZa=d_]RU_O[]>CZ_38>Y]RD\OW.EC88D1/TDf?FBed
^F>8dUQdd-Y(EXEN0_X&6d=UaYU+98WabVQEdQf0fGI/E,d_gF3:dU>9<Z_;_35Y
IM/YETC9^P,LYX<Af92IBDQE?I:#4/S/fd3+7]a.]V2_Gde.0=?)Ac81CVQ>dX(F
aeGI1&/M[[X;9HX&ES=V3bD89gPSBWa+O(O^:/eZ.])MDgSXU11=J^gX[Z[N([_N
AeF,,/d(ZGWbT78AXN3QW2H.@XXG#U<WLP69(BNFYF/RJ&F0>,9>E3YHTLH7BZB)
C/=V;c&>Jc?E8C@L+@W55C1IRH:D\d&W59BAHL@+\?>^S)QDaQ2IYX_Db.T3E@S@
(U[3+B1S-&eSH+3V3TQV,XIgP)L@2A>]ffKR>JNJ2:c5E6P+7(g1D0e0dTHHaA2/
MSDbN6=dWC_e?MN0-?+=(-Z&\BD[B[LMe;<:#39/f(.ZIaAcU6E(ULZfAMR98O<=
c47C5OHaEbOF7L&<E?2\/V:D;,8\FG-VW(f8<C.EO;I2b939L=9dC+OZ:fC1WA=Q
^&:7-,\0=>gH\1(\cV;ce=QJT/?&6:c8G3]DEQ7^KUg&OMRc_E+F&8Y2f)f&(=N#
N-.<T670T[\/Q++Q8-].W:Q4AM36(MZ2;K#QQ@&56T8GGI=[X4P8XU37b^aR.Ufb
MGf=9WCT\0U\f4Ae_#SRcAFN@,V4PE>C7X=PQ6d;FT5X1C=K#7]\W[A[I&=JbX4@
5HVEfa1L@eYHee]SaOda>(PM2=D)EJ)486HJNdB^Y(4M66K#7]dT2CB>AJB-657&
8YT/HF@B=Q=BZG84YK[:+VFC4b)R-eZfDU8b]KQSV#8?8T2;dIMDD[Y#dZO.YB3g
&NS..aY(:TAOcH2X/C&RO>N_fC)FW)eSa9H6?ZSB422G&47QXGL.Z)cO_/aQRP]L
L(KI/gLfY:#S-9@V_4g-ac#DNJ3MWA\X#;8]6gQ-5=KGQPC]Q,fP<PLS8;_@^-MQ
4W7/GN_>&X(f/I;g8Hc3VcL\ZcDU,4G3:[912WfPMOJaI5dN@Ma9.adDSe?VX3+:
\^MN3fd?g-]CA>?\FH?MZ5S-A&N]ZMTOYM77Ma_PSad6IJ>XYMd@bH#?ILCXY]G?
]N-#8-G#V=9RaC)SE&PYc>];WAMgCJQN(<[Q](:8_FVaUI&O9(Y@Fd(3e]DFIFZ]
F=#C;X,\Mb<(g0G+3(gN_]SEVA;<8Yg<2.+QNI;TP+Y=6/C-GX0Oab/7F/VBAdM_
&NR?dE_1F<:)]b,5Bd6C8W1+MY58&;BNK]X1T+#e6DZM8a&DASV[.J=/GE]gL#TC
Z;WeZ#^-1K<OIb/1-9-\@3)a7O>a5?C1_9JKZHC8,KY:R>cbI/GP)Y(ENd:J=\QL
XHJ7b0+bUQT]+:/NE9O/73aZ^-ZIV,EWMY_<IZe?S@CH@NAdcR:R.ZT;f@EV.9e6
0_=BeL1G04ZDa@T..;NQMTA20BE/0Wb7&Sd9NN[KRC>1URB3NA3T+,)Nc(Y(60M+
ZKPcN1,<c4T,^B6#HP=Wa3AV15MT:W8:9]BL6#E6dW<G5Ge&;=#:G0f&4A4WFaK(
/Bc1#X]RMHRf&@57O3VeMDAPf051U]#\[KLQ.e>73>^;@TQ6@0,bYAHAUFA7-D6;
K<7f\Z2F_[A[+/>ZVT#\a\K(baD:HKORH>GB+B.<XY0[H<A?:13-UbXE7U:FdIgO
U1fa)MGZQHe1U68<1-g=7Z4_LB^6\^]g2Y;2[dDd]QC1-([,J+8B(GMG-4KI\.:f
eRK)3A7SQ)#>6_)8S+d-#5U(7]-D<bO<L-&_F;/A+KJWf=V(be^]YJTd@eK2-H<R
=&U@])2NW>:KA)6<&;5&g;>5KaK+e4)d6b,9[JZJ>14H#Kbd3=D.7K3LVb)VPTec
HK&fWBf>B27<eU1+.P=IVAMBCY40RI_/I&CZdY+bU<E=HKO\EOYP.J4Z>O<(#X\@
W7?R[6fKD?U[9AL^3S+M+D?g3&44I+PWAN0^L^J;aG+BE,4dg)3F)1L[GGe-@IJ,
W+?c?R#FJ,K]MO&SQI<ABH\[12/4,AE8e.0YGV<<+>4;OfYUWbKXMM9b@f+G5SZ+
:\+E/(B/(XUf1eQTY)V,c5_AG]?a9CgX^EQ4]e1LRSHG[Sg5&b:Pg=KW,=(S.#<.
C9AI#<ANMOI>;?P,cJ]RM&TG6Wb5QaaeWN.+L[_:@?EYG=]gV7S6N171M+VPF.e?
</-&3-J8OU8GF,\fIY\,X\a=5WC1SN@Hg<b&HI1G.DUHcRW7EY[+eY-bGX71.-Hc
LcPW2KRL\>6dgPISbQ,9;2F)SeMV[;K300,f)>=XcfKL.Eb0bTZJT1]X7U6X^_^^
-@TQ^MITa,F])T.BfAV#^N418=<2#G>XI>AO]V;fQOMA?A(J5;YaC:LfIQV36f.a
7G=dBQ,(RONCa)283.YE\4Q(aXE:eJ<IV4)Y[D]E&?a;XHCVEeL3+^=4La>=573J
H,^GGMYc=&</;\FD8L?G-UUF=>>f)]QT^>:=Ze<3PAX06NL,@YDfg&V3\cW6MJ,O
X8BSICLULG21Tg;602@.<#c(FL)S8^++.=P0B?)T45ZP(@8#de5)2=5[]JCfF+@S
^7KbebHY:4[(#T]\UA@f@V6d=:a]g#K(7M&P<\QfS17/_P+LQ/Ece_JS[XO&VD@^
W&7(5SU:I6Cd=9=eK,M3TW\40EcQT-BR@aQI>59G^IdcbAbRXKe&IWF=QS5X,]U6
].TVW:A-GKDP2?K4<c6bF72c(@??&g.bOHW>=+LBCfC:V5]g27[RC,A][,HW4T>Y
QXcZFQMV3J]_TTeb9IZ>9SS+6&V(e<7YeLLX(bQF-[WA-_(,+.M2G:J&dKcR6K\F
g:2\Z[7UYXY6AfaLKYc56N<S8@,eN<J=)@4YLDUM-4e1+1O6__DWJ1OffF:G\.[g
40=<8::36A:3QM\?+XQC@H.4M)>7.\g/6-J8PKHTE/]XCQ?JL--c=>H(&[CFZ0QT
2-&4SA^4Jg(DS&CbT;b:)Le6R6C&-8HEcH=1,6<?7b5I-?WfUZ/>.UTd>I8DaXL?
/7Ja_C/<(Z5bS>A,#Y//Zd.I/1:K@\b1DIDWdLM=&^43)58aIgabGTZQ5M3d)77>
K)\W41=I2XGgGW5<9FgO_-:46B8<.&&73a6R(,G,2Y-^V8IS6_5:\03EHfL9a]2J
^?VZ0YT,C\ObMcYM=S((\YH391>a7XVBY)XcYb+J8)1eNGcTTeKg>PV;IGb.f3-S
]B)W(;Y/3:JN<?-K64ca#OALO[FYD&8YbOC@..X/AP-V+5Sf#KUTOQE:6;bKd=J1
LC#YH.;e#9aaM#b#=:GG]YG5\Y(266HHN3Ic+18cHBZL9;AP#H5P;P7#0331AH@<
,TQFZd\[/S62fT4W@>YeW_XWE1)Ne@F_>[ZH\-1JQ0D1YCgVHDVHcQ_f:,PX\K0E
0-SR5M8bC(@:7U2/[.7([6I]CSaOg.)Y@9JJ@If.:Q1&S@#9;(F?:/Y_[.W-531J
/\JYZ#Z;2+,fCB8Y.@Q/A[ZeBJ3g+g,XFc0TeO\C7X6@=D09+=7-Q.CI1c7/JVg#
E+59M-U\[ZL/I;J]42](>I</,<MQ3f+RI&F_WAL]:fKKJ+RO_5cG,9FFL#g9BTY\
+d7J,2Sc+Y_TV;:#cbf>9Q,X&b_;IgcGC#H7df@BLbb8BSJ?&>DV0#^32QJI(GE0
&K3b;_]6Lbd\;7&+7RZXH?&FM>EB65Qb3/MUXK9.]?.bc:#PW2UE^?.R83]/+Hc8
=[A76#XIV@;a#fJG1Za)4XKRVY:Hf()N+R=gJ4BI1/4:@DU8?;E;aSOQfZa&L.M=
F_E_)g&EBU8W9YccJQI0b_TfX0Qg333WEMS;^.@=XgP31^>?A_-UINZ49OR#(0U;
)JC6M(LLA3Q:(,;UcU[#feXBJ]S#)A^caYc;-d[XSd,@ZHb8?HN^M8J,BOFgJ0DR
S1e1B1VD&&_d,cIYcb^2Ue?EVPGVT)EL\W?aX7b1F+66IUcO#WE()BJHNe)b3G0Q
(Qd^7=IM,R^6\Q3Cb^UcJ9K4e9Qdf&1O5]W\>]H@=@S)8Z64eU..J5FR\MR\=)OJ
dg12<WZZ48S3WKT4<.V71?geYCN4W\WZTPU):a7gdS/;^g90YPED=GEDOS\<B@K_
Wb\TD6d_)CUD#Q/WfKfg0\UG6)]3faJ)/)7b[(_X^L+W-V]7d1U<:G\=1IZ&;YR_
T3/@T=TFB-09X.JbcPW&Q@Z._C][RMJcg:\BA(OTWd3aVRM6SD4V9XaX<_+,9-1V
5e9I<K,XUZd.3>#@H]9VP(P+?I@+AR-\Ta,):T)86_TJe9MPS=]G[SY>:RAID2&b
gG=0MAQ1bc6CRKE/5:1(M>0MA<&)#::A9[:(A+IK4.K(dg10K9LGa\AJHYf>HIU\
5=6;f@&EJaTP))2+Z;@3[5R<LV4)H?[eLg,@II9^&@8F2A6?#MBTU_H+6K6dA,C3
:a)f7K=[Ycc8Jac]JNYR6(WGG@^H:@]R#de,O2BYB>DgK)WA^f9&aYX9f=Z)=eJ-
M(O\Ig58?8c)G-ebV9/\7][809S]S(PbY60GGRIgAg3L[;2QCIT:HLU9(Z-C/KFQ
@Yd23Lg]O#1L0I7e3BeK?b^VH/1bL7F]8-H[XLKD1UV15?cbE[\NaEG>QN93e@Dg
6&.H/DF(-RICPGRR-58^-F:bc?FQO24E86_.XT94P9K.5W?V>W,[U^.f4KVDB+&V
)?S9;9?.)R-NEKT/XH.V3]7IJcK0eaaE);fc[L>;OCQ8SI(IZ]_T+a#?JT:G1/Q\
QI(]>@Me.MXHcDKf(G9H:EME,:H6T5_G9U<AObN8,fDQKH)8:dEZA6,O.EE&O<dG
-PB[8(W1fLKPG.3,TX00Y+d3fZC_P2OH)eD[fD4f9NPUI\QID-G/;P@Rb)1L^84F
/Bg42ab@fI73/Wg:4>(E2:0;SUaFGQGIgAT+Z7.Y_d4WNC:Te5LC#RU6=f8Z1IOZ
/d&EQ>R9VXf-Z^,LZJA+,bF618[,K\P?0H7?J0_X]O-&4b2RTT4+,,NeA<S-.If0
?SDU>M)3Ge++8R9a\;dL7g.B+\b<^^aS2c=,?LYYc+^#JV4CL2bJ&2NF?LD7M=VD
=De@[0e>fU?)_A.Q.c_^XIOC8TaH)M4g0Hc4AL1=<8[Uc]:7&#FQJI3DL\IDW)\4
\,bM_]W<>9-?B\0V6>__fNQID.8E,a1L2SCM11_4-\fTPG#0R/4Hb-/Zf[A(bC^]
LCG7HeUIO1L@g1#WG,Ne>_MYBX;WJV)W57=b;L.,/C;1a:3+2GOe9[GV_S/KG<11
c&^YBX>M.(N11.c/TE\GF@=O@2>Eg^ag_@=>c:@=&)c7S9AI2Y?I4/L3f)4FZbX.
WHb<>d18g5YV>g&?E-C\<XK607ZI31bbOJM-HX0L47,@HF0>FGdbMX9,^OB,L?()
OR5^PCMB03P)D(?-QZB@\;HQd0\?KSd])]F[A#X8RBNW_Mbbgb=YW=eF&3SN(XF#
:+U:b?<ZOR&fD?YOcS2C?KIPdCDJ(R\C63BG.7G.8b2=LJ/,:da;.^0Y=92Kb2/]
]<5.:FG:PB(K8CD5XH>NJYMAcX5>YEFU-fB>#fa7Q5=F[)0K^C(,^>?)LRDd+g1-
R5H9N;(eGB)WZZ9=HXLO4:L+:ZbH_Q8Cf_&^_?.E+SC^/YYK)J.[1:\LLcBR=<_M
62Z6VD_V2REEF]H:3)08d6+Kg6\&SE<]G4e1eTK2Na)(,<_bZ.S[VVcZJJVJF3.3
.L3/LD&@MR7#F,A9]DF>;JI(;W9LY\HVf52TV=UY7J2GN1H1c0[W,-HA),4GO.5^
O#e1_5CPSS<EY:LL;e9KT4@6S&FR^61BLB=ME=J\^XJU6X7^4@EA=W,?V(TDN2)Y
fWGFD0H&5/<#RL8fZ:WG(^KMB40[@dK,:NWQT1Z;I>:e]dXbNZW-35=?XS-dM3-]
JVTP:AW+HS&A.B_Pd2K8N6PU\/7@IN=]=>)EeM\@TXFW3+67/^d6LHVR,5@EEN_F
279W6Y7RaUHYc3WCXYO>d>4_fBW->/fABU6:UC-?VQ=HA6f0>1DI=6Q)AbRLf0\6
P;_0,f#LL-QA>g<X]D?QdAP(39@VPd^eDY)J90.&KEe-bcg#@7:_TL.Xbd[?J]PO
7A5?FC@K]0QcDJX)\[BX6,EIC5-cL=1R.BWV[WSKE,cB7)O5.<-Wd@[)H4(fJCIG
AH+\\1E5/3L@IX-0+27b=LLKW60ZX,Y=4R)+&dB&TOW>c,cS:FCg&R/0=2g806#E
RbC@gO[Z6g5eHT:DR8ffLbG+cbQ7=>T#S,SUWRg>=J5/7H<YX/RO7G;:eAL;0CUA
cQ[D.8W6VddL[gdEc)8XQ\W?>3C,WgBR:?#>BKFLF[8)XQaS]I6(eD7/,.(:O#MD
IPMBD>;,[YU\1A9b)M4DCK;WB\?O-(>0B;e^SB\JPbT&35-AgdI7UO3^OcdFA2Q+
=\5/\VOX7&459I#1I?_#bABU2[.QP=_XC@60af]a,Ub:9>KLc7RGGN8U)Z]<7I;1
,,-5B=^5:RBZMHTQ<f+33JReGMLJW9L@Z.S>8L5a=S/<CV;XdC)ST0f&O\6RSG-_
,efSX?K@,L1]4@AU#FHM?<S<OcPPD;Q&C38HbQ-KQXPDK@/Q[MU(T3BF&H_-96(R
>FC>AbI-\W/#g,5#>.U:RR)Mea[RZMJd5+0a:950O+P\;YXcB=V0E]:_.fO>)4D0
9GB6S(Wc0^FW56B(.,LNgb(G.fHCPBC2/@1c3.[a=G-Y8,@CN5VdA@AbaHU?2J4,
<V\+(D9/.cK6.0A11?_3[JfI>PQLNTF\HZABeKG2O0SWT0X9@V_Kaf(L=U<B&UaC
3Ic+@@4JHQd1T#HG/+XR&,T^DCPVFEUP397C&;JJ;J:NS5;ZN):0Z+F(a54^d+0=
&DMNb//;c_PG#-BGdN&+<&0^_1E0@IbCW9YTa?XPAP=1fZ9F6[O3OMP8&,gN]:]M
Q[N<LLI(L3:^Q?9C(5NC?/&WB,/L]]8N,8,KI:P>R;4Qa:De9?d(\Y#R-e8):)eT
VGaG_B9XaVIC77Oe7;[KMg-]YK4?499]ZKd<YZH163Bc?RMgAQb--Hc+OLgO3NQM
:[^C67::OSf>?T1IfJ6I^U(B5SC)X59X,=QBRXacWJ(6E9RXbVX7L]>f1b-:DP6c
+()G7VNgDE.6;?3-Ja85+[U,=M/8,P5:(VGINbK,95X>.S?fg<Hbg(;@d>>Y]BZE
.cNdZ-R9I9-3GU7LUP2E1A@92T>P--bW8afX\.VFM^D?:8&B-5KXQ3&fWQcAM[<T
TSKXM_C/VXdUX?UKDHWdBNOR]&1+<0(CT9We-F08L+;-VK1X;IT.4G,+0Ma=WRFG
Z71D>9-8XOGZKGWZVZ;f[N0]g6^+1OH@_+A=>Tf,^>O/81??CP,+9/P)@7MgAB-b
2_@1OFG@K]/RaP?</1_P34M,04HeNNK;Wg>#aO2K?&2]=79(eYfH2&AMA?DW;d4M
L.E()HHD6QYUA#]\fKATZWeF_E1\#LcOX996D<)#,7+35dcaDd>(:IdQ5)Ta9JY/
FXL5RY)_NL[e;DIZ4XZH+C3?]QIW[6K5=(&K9L9;L\/OH,?IMVN(R?(H?&9<)HQ<
IS&TM<F,MP?>C]Fgg?E]:1?RLZg=V.-R3f./dN;XA@aGf&3YZA@V0Te\_fTa1UIS
,I.;O-+AU+J:OI?3D]=fPC1UeRIVRD_bN/.N0>0BS<RK\FO]e<OY1?S3FQ60K.SL
L/;Be.G3G6YK]PTWZD(\J/HEM9cAH5\DOa6_[Ea86gf+,WcHLY:]H):We9+YKO;\
_8R_2ETX;aK@A=#bO:LCE5N6@6Kg9>1(Xb+8D:a>()8,3Y57MS@-;NK:+H+;]aUS
&[55\=4\:S)0#@@3D-=5]NTO2@V;..(.@][AJNPO=\ZKO3WLf5?U29X@fGd.6cDE
_;I9SU)?bJMd>5gB&^(CL]@#VI5XT>J)(P4e3=<UPI_<f+HXO@RNJD[^>N,=+Od8
Y,,Y9^E5/K?.,NR>=0/,-adCC]3,\.^^\4.HG\MYG]g8]&YA><VM(?\Y@bUS;d,,
#8(LMND,+H^OBD[23Q=N++44UAb/)T;8L]&e9A-C[[]L-Q+A>CfZ+.;F=8,NM6SS
A66V2fgB\EK3eUP<8@23+0CG63b/]O\;JLN)KQBX]HNQTIT#gG#g2gPHf5@A4b4[
WIJ?LV6Ue[+&)M6=70)EX#[/_A5Z,Y#)E](:T&&+6\,VFXQH)5)6dBW+@<=c^3I2
U41,L)R)0ME)dWHQ=Z#E<CE3M=)2@5PZ/8VG-UXV/@bA95OJ_QYX_+e7-U2O-FY:
HIOLF)SUa,Z0E9^8&H81)HQ,)AJ7Y24<R&8d.]LR#V(@[6bY&&<g.RSKK2-O:=81
2<=D(2\4--(a35#I9V;QJ,[E,FLC]b&]=bRY:37B-^TMA.?@HMU/6L=#9LJ<fHb?
f6gReaBdbK_;YTC:DHJ^,QHHC,.6,ZZT)UKZPH/++Za=[GZM.2W&@c8JLJ<]F1F;
9^M<aWN\F;SX@@5I43(aK>H42DC;Q>7][@--/;3Z^M)W4C0a:H/1.V2g5M+9.e13
MRIR^_5;4:RNC0H][D-6MI3EYYBG<f8E:(_7;Y[[:Pg2B11aTgM.XG^E[a-(FCWZ
&&&J>D(X7Ac2g?eeL.C(0AU]0Qg)BWLI#a-1MFa1E]TM6>=\8Z78/MWB[e;S0T#P
]11?F0QEMcT@\>-Zf8eRgN81;U&,_2^Q81Y?G]_4,KY8^=]d@6Hc<)25X&OI&;QJ
6-/Y.I[<I\-/b/S#[A4:QMKY)-aMTYQd=7JDM]97bOO40ABIOB2XfcJCA<:(^;@/
W4&=:/>)LaM[>e?V,BQaCTM:9JT>03VGc5\)WT&BI@Yc,deE/B;O8V6B79P04K4Z
[:O2FUL&6JM&KT+YCbCIHK:L6^aS&]cT1K=;g;GAU?X[PW-_9>?XMUPV2&9ZU>#3
0?1KG6?MQ)+H;f/I5[g(XVP)LY2TWfO])72?VI_R1HZLT+])29N>8CEdSL\N#]&P
=Z&>>KX(JQQ>-b8#,)ES1Yg^OYJ@6/+[]VV.R+]9:,5>5@9=c:+KeHY29&<\M\S)
#-[]MHbCA,Z#OfN;WS-)N\B]\<Uc1=5d-EC@9\TO,8GK_+EcCDe7AVM&Q4HGJ4a=
eU=eJcc/TS@&>P^.8.:3FTYB1A^O/&SI^HG57>1b,D?XA@#4DFeJ9NMQ9]GTTX82
TVM)AN__4NB7MeFIQ+,A#XQ]eDU=<KR^I:D^gEOeB+8=S6F,=;D]FS4e4#\P2+D?
GEX_^EU.WP&-LSbg/)ZC\O8T_bX)4g:/7H_f3#[DE#8Qb]<>T4:9XU?[F5L6_)bN
I1UK^_B&0P68T>SVR7C_cA<:V&38,1\J#DSKIE,61dS^;2W^/OT/7&R=.5>.ceLD
fUCD@<g^:/GdU#Z[c=<BVR<J6#;_C;:?B8HHG?EO@GHDORLg]<J@6^V-Qd:;;7F8
a@T^Z7O9:6PENZX&P2aKWLgAgSVBe5=Z0^U=DS88LN2(A_72)YZOPDSO&3KEb/JT
D_cYcN^^0D1N\;UB_);,W)W-A;4NJK@>AEb:@O/<_O>7#\;@^bbdd]?<:7\U67(P
ALAd&Yc4LU4?UPTRFLTf13gQ]S.7.T^56HV0:5G/5_T_Y;^<U#<aN]V-RMJMU6LC
=##&0DANaR,=\MJPME?)g3CZdTaSa#dQ0SJ-?YU=Qc)EC9bb]WR12S68+5B+XU=S
RAP9?/4?,1O-;APUc5YR1Nc[65R21\84#.#)5.f8#2e4+0[^;2E[-/M.=gQOZTCa
Pe<COEP69.]6Df.@IH[D:H\+X>f[MD;a\MM19BCQX3H1NAH7FTM(gL9:-FMD),/6
\4R@I8eXO<AGFad4:VWf.(H)GY0VO:U.BAB9C5)gR1Y>\SW[e01e>^Fa/,2YZ1.2
+fdWVfG56#MX>^0GI_(9UIc/gLMKW1O(e=HKNaCa3-c&)?=<VCc8P#ebW4>L_G2,
VD6J)6838OWSY[5<Y8a))R/<+fd7=V#Hc?ge>4A+>WLPDX&_Qde<,_05Z]e3DXY)
485G^CR7=;gTZO<A55f:_M\D66I@Jd5^67RNN-@05FL@>7MUgg(7\4CKU-)6dD)T
&9c(7U/3#NOK5I/Tg9B6BB#4:=TGfe\_bgQ&A1QVaRAQ;4Tc-3<N&MKCT:7<HZRe
]:bR,_68&FDf1A30eaPO/@QB\[FdH#Eb4M0[:Q[+fCfOag@:-8SdYK0gX(7OG242
48U?egWbNdV]A#YLVLJ&?:K?QG6@JK;VFeH6KXO(2)?&F687:419g.ATI/3PWAI)
7.?a#J==3&WcFd[>:,W7XPYQ:\.WQ<:b:-0Af3.4)QDQD-FQ8_g=G[Mb&U:aSMB.
7dZB0:_)d8f3I-WgR6P_MW)<@^]7@eYW1]M)+@]&c#/\J?EAX\C39(6^S2LecL]a
ed#:KWZI=TO[5L>6a^_7.\ZPCR5P07O=fLBVX/15Q^:M2J>O-/(cJ+M]8^K7;;RK
5@.85:_)K8:(^T&;3SLf)U&OC3Ka:cb&N6Q81f]PbSSVN;Y/ZB0D5IJCNL+8OQg)
]__6C_S/\UU?N_-NFg#5L(\:7O^,XZ\<44C5XI&6QP=?1SV]KQ+H:O\:5DIO4)VV
;H/P;:RH6L6T70)<>TBUPb/&bAb@ZTO&0]+gg2L:5.e.R2Y3=&GM>W9Mea97WX7?
-c\;T2<=LR&L.<78bgP5b9U752?fF>IZb9P23H-D]F<X\_ecFJ].(V1^f0->Y,.+
OZSfSLZ2BEXB5X;Mc1.8g4RIB1[._W5H2&2C79<I9Pf).F/A#-73_CL1L:0QNfJ/
@B_WgY0#3KZQ<S79(D:I=M2<fQ#)7H,gcII&/c)T^D]f410DGfS1X^J0HK[-0Qf+
cgGV3TXQKGXQ<M23Z&V0;,K2)HA;,PgBX#[0/-[V_5IHC:C2:M5\PGWQN&K6=d-A
_1JFCZ0S_/.#RC8GU-0_MCB?VGCN-1=L?YRU\DUJX#MM.#4S#f[QgfK10AUd3E4B
#;7;6;5J7<SMKNQEE\<]+&c+C8]e;dga7Pd\PF53XX4#9L-N[7Y<HR>XT^\=ObZ5
<CBf:(0PKB<=_L<aOWPSbRND,.#X@1V,g78TNS53A[SCMGb7N)P^XU2=-UC=gg;B
[/3FM[-@SceOQMgg9,LMXfSK>\43@4c/GIEI_PE9gQY.Y(fV]Y1a##?I20Q(Y,@9
9f((H;Tb=<;XcBF]SHC;OK+#Lggf9B,INQX-[RG81JLD8HAF[d6>-^,-BR2?A,<a
<:..X\^L#H#C+6<IE>6#5D:^#Ad2WD+J:-TA5d;Vd]>)[^AOg&0Q.Yb87KH@(J[]
c@[RKdPH]Y2)IaWVUBF(=4CQaB.8ETB.C>SJ>R5bF,[(:@_A<8G<.LTX&Q)c?8^#
MJ0]6?F]<#FcNPW@ZOUH&GQ(H#OZX][RAA>_\f\?O-SLI;cF4<Uabc/#^ea,]R7B
ILb/A1ZEMT(V,Ye)IDH@WcF:7HDZOaOU[gW8LAeA8UR,;35DeVLL/?N=6D_(f?VC
+dgg.,),_\H+R/bcQ:H-8.5<;Y\,gE[fT/)#63IDDg07f#a@4ER.39.-&_ce\OCO
#LW6/6Pd,RfeK-^2&NF?]beYE]3,7S<e)BBULL.<3-Y8)SK>&J8Eg9SP087-K/bP
MCKW>5ECJA@7@F,#Q0-QaJA\N#_Z4O_?c[15PN;_ZA39]WTXNg7Ea8D27,aE[ARD
I4>)Y:eFcGABX#?,0.=?<YYK)91ZVKb8(+K5DV4c,3P?JSF\X:AD/W<9O(N=6f+6
e2CZ00WRU8Z^ca=5/#B#H,J^;((#^/&9GU#:ICH?Z4,gGf)=[R._,5fC8A]=RL/R
])d7[4+&a@#G67&0627VV;IY>_;:P5A8L?[5<B.9^e])gGPfX14=93<@FW,?4&/Z
63I&VK?FHUH-]CcHFA>7J5U4aC=QG6N@ZE?+BMdUKC:A<\5/&fZ?6H3CUR0FHW?S
T;.d)E47E;O;781:,,QQ5<ADNED9>7,O^XNKCG^f9-bI,[db1A,NRY<gOdEa3a=&
cY5L<eDa4A7C>\YW^c<39e<;@a&Dg#2#SRUZ34aedaQb2#GJ>.31[Z/.?X^F5^W3
#+)(15d[(:Z9&RVA]P>Y=V=3L@&,+fOC>S/c&K/J(&L#Y>?<0:OM-DK58M.CGER3
Zc]bWFJ^X3LS5bU48NLXS0WR3Q(V?_&SAda=Xc]5WfEaSCaMe;VUH@<=aK+e\:>9
UEV=Q@eJZ[YHA[TTNe1e;(749_S)2T:/(6B.@fEY8[[ARJQW?G]Ne4??D3JN?8Vg
e0eHbU(M#GG0.K/Q)Sg<a7W?G(@(@:.fM#YJNG#ce3,<5d(QYdcFJ0b/0G>DIPIA
f<GI>)7>Qa[,N[Ze@e(&5;8RPQCUA^C_+TM,0GTN^P4\4:?[Fa4/S8=G(EBR>T;B
3Lg>_R4HLIf:FS#+.gLfC,DF5g^DAN>__C?:U[c=HU1]bLd6+KY4.7Y]Q=f5dX72
S(]^Od1f+[gM<:#bUSUbGdeT64fA7OJATDY(GB<MN).42+=0<X&R,3T?Ra_bG1.8
YNQ4<@C8d\ZF&Z9=.58UDd.<CQgXC8ZDb;<(-b0?^ALTfg3S4??7O8<A0GVd#BS(
\HT]PJTaE66]]C0\C9/D#/D9>91,9X^=e?EU6VeSUb#;@Wb([K7;VSO<5RT-E&gU
0:39Ge.79U()dX#3=Mg:,7TC@RY+c..E4AK8>Z3NIK_E3L_b>&K+MW#/_/=e7+I(
McM8YS72=I.C8;X67Q7_e)86GXJ[d3LCD#ZcCMCcEQ1HF8/(]65+<26L20dPg:?c
\SS@&@1T<A-FC&ZN+HX\/TFC?gWT50SM+UIG0M>BbDDGbc_85N5>d5g;--.QGL1F
JdEL#?)ZYbQ\IKXQG[4DS@XAF\PAH3CHPHDA^<S97Q>e<BUX7a&A5(V:#47XSJ.H
>aZLCZGWBSZ#[>Y0N?G2Tf+9I]/NI+M),Y6]_Ze7aQ0bYWd-=0E7-C:OC>SfI<9>
[0HUI=LM:B43C@A<)&LO50/^@GaNF(-L1:=&a6)8IH+6W4(97)+GH0PfYfOYWMM;
=\,[BU=R]8UDVg[4_dGCX.XacY[)+5aWD0+QV]<T0d)E2g3?EEKD7]L22cIB?b?8
I=IAECB+6^;OPf8b.([3?E:?<a0aZeLgX^ec#a,BQ&+#G0?^a,Q;KV4g(d]g/G&c
9J=WJg81d6ZLPa>9(7-PAabSUSS-N:EC55]H.;gZI-b;I=#PVR[/SVD@H/Yf]\f6
2)adcVdTAU18AN6GALZ]A2]16,Q6IVSQ6QGaMX8#bO__W>^IZJ+a\gVU?>D&9X<Z
+TZHaLF1@[aYLg2;F5:I>MUIaQ//7,4?0cFF1@TKFW<<?2+@Nd(JJe)JZ)A=]#\8
YQbBP4\9ff1J3O>RKTN^A&/#O<.bK-[U,-Dd=bL8-bS-GC6W?9,gX-CI8H_[;FBd
SLg3E2864(NKK+[Bg?0R98HQ?FfM1.#Z\bDB:LQ2W0aI-0)1)cP3KK[?\WH+6,Na
^_b0d)UbYKE7.]2J>:JG^Q-BS=:cX<fH4VL?ZG=1G3+W8Y6@EXO4>/,Jf^>0MCA.
&A9/Q3?;S1<;7U4R-e;M;24\\M^MDdT\#2VLS]T^L-GN>g>@6>J>U#^PDVN@H4O]
P:X@\+YI:QO]]1NK+:0_(:eW:e4NWIHf,aL(.6@GRPDFFT&)F_e#N+#Z,U,:?^E-
,89A?)HS:2++U&g9LfcSLc98aIYU#5VJ[-ScDZKD7X/XX?3DE+C/V<OcTCFADVCc
[aW>g[W[SeA^.F?R#fN4W>R=,&AI:a2+J:bRN+bC>bVUPZTgg;)UL=)3.bDb+PWU
&QIZ57bJGZDWEf&X/5d,E)QbbBC,?7Pae:PW_A[1FdMVNTK2(W#8YWg^P/V/7^D1
B(-9>^:_\TM#>?S9-ZND2YM/2P4dH3/)VUIYc,9aAIB:bHX?gT?Z492-@<FJW,0N
IC/SNT4V?UULF<VQ5E7K-H2:ZRRR.+,06-50J=eTVO^VM,Y(T&^4A<<Cd;;]0K(<
cCLf0:.GbeZ)_c-4V>T0N4A_bO=./3KL46])#9R,24O5+=NI@SK[<P97,@)]H2;)
U#>\[WLQ3@Y]9TR#(37XVG(]2eI6_N#/3DH6IT43XfLGecXN]S_]S1&FSJ=I)CcU
0)D>Hf;10IJd3.VdVdDbN1DPIGGECBKZe-Q[=Ig;-;\3ZcVdHN-2-C()-T3M/\QQ
1MQ(9Wc]D.<cJ+W#<KA\bbXRfN)Z^CV].B;&>(=7\9)5Fc5gde&2^&H4BP&?=KbN
ZVA<Q^II_=R7/)4D&9:@edA(KD#/^N,2e:c9c=[R2Ac;&AIORAFfa+T;5F.b01:7
WID9BcZ997c/^K8<=IEH>N;_1K:28RK:6GA=/4>L=K^DF_0_WQ#WX41)(S4,ZGM7
-]7O.15[T1Q5U<AR#\42g\B3Xd8C/G\F1,(W+XeU&fMYWN&+eb;])>ZL^=PAX-K6
1f/;9d>]8c07AZ,DB/f:@&KO?/V3:0(\/A7=Q883Q51EI\e<QfJOEVGCbL/IU&gX
OG+(ddH(7<G<=S1Z1HfBd42QH,K8X6::0NV:<=SfHJbSY>d,XVeO;Z40V?7&@9@P
)]WBWO[b>9Z-RSVJ=H[^;)MZV6GaN(L@X9^UN/^,_EHC1S3Ob3H2/D5[#bT(8G>(
Bb44NJGEIDbD@TE@H?KTGT3dAPC7FD^cDQB40D8R9HZB#?>F>6[cGNf]09f5MYG7
YWJ:g&SJ1bH9WJ.F6M97a9T6-,7XTELEF23<M4E?QTOC]]gQ831GN=@0=PBd=Y9\
C?F6GSeC@Ab@ENIEHK4AP4X&8E61]=[BVYEdUK^Z>[^ORZCJ+Y=ZWVaF?27EF-NO
.60DTdRYL5=3S.Z-CY\=D9g;d[d[QX/dObIC=#b(aW/.>Q<13):aS+_O_BeL>Y>]
#LKW=-3b(<8:Ob1X;IFgH(#KB1f@IJE7:@W]3]K(cL_6[N@A6.^#-1QVCb>\d&aR
?75a2<#N@R3[bQ:)dWDb]31B]-Y?QbUc]\>9@]#0C_]4aT,+I>7(?L#<M10@.+@L
R&Ob(fF:+DN8O,2XHMP[b0c1SfCd#_ZNd2H)MQQ?KMD;=/2RNQBE^1:[LJXdEdU2
[XYedHVW0;>HVaH2NF@7TF#RaD@05bLORegP>1fM25PXe:XI8V13_13BC5XR^ZGa
UgCTMX/3.]7YdF]R1#FSQLW@GL=:6Z+)F8aF5fIB+f=J3A<.I:[)_<=0_IEJ=30K
Y^WT\K<#\>RY555J+3Kf\YG;Nd#bA++MADOa6a+6\F)a_\1^c_BT,7#\Gf.UN=R/
8J^8(@HPB1RFK=KHOVb7?I[&:e[aKJFNO9FITZRdQ)1_&N?X73+1\4fI39_OYK,\
[Y6,JVJ&4D/^g)N\KdQB8cPg?(F<DQM@/G@#QEE),WMbC[]H7De#[63d-gJPHe+a
N+6[&VPJb>Ad?E[P<,K<0JXN7B2d[UUZaG.;N#([5K,<@^&3#2P7]\(.J;IL,H01
MK\Q-eU^@=DMZ9O+A+2;f5,OFC0=JAU3[\UKPc3eFYRQ^#_&-K]AeH4J.45PecA^
ISCP>LcKeIIGb^cE-.ES+IKZ8f&6@0DONcf_aDQF,D(X0(=^<^EXR0@]e3>V-L[Z
CReS?IF.]I+TN;.&6C4b_R#C<E#/;-U/-(#,[PWg]5V&)eNF4>YJ(ZU.&bNUM=TN
^=J356\dY=VY5H[]5:gX\T88X:.UeNHZJ-,?9IfO-F.\18N#5dR/b+eMJ?1gS70U
P#(UaYCJHXQ(O30D20JU17J=R+](NPGUUf^#O.KU=K:,[VR<2:/5,Q(JDY0(63<F
>.#EGI4N.-dGN7N#?DZ-QZg_@.01X0NcbOCK?Wbg]VeI&YRY^_2^c4)aBQ=(R</?
[#QD\RF(((=14GS1>NT5L@(aR8^2TQ0#TY&U1fJQ\Ve][,:TY&&La/^+1,g08^@L
LG9>aJ5AG,[^:Q5H(7Rf9d/?AVNW?@g4&VQCRC#)8:9]:A8;LP-N8ZXT@CT6IH-B
c?UN6S@JPOH]_cN.F\[f]_?/agbaU/S5HP:\SU9Q2Z:ZZcVD1QFK^^EfP8XYUG<5
5c@,B1SI[RPW,Q@PZ5CF,B4@LVMYR9cge^UIO]a64/7FV@;fF.K<D[U,@e.3g-5K
XIYZF(R3L@dg/fB;[SU)5BC\,bS8M]U9VSCSM\^.O7JgJIWFfV73.MCY4H3R[NT+
TMU7bc@Y[K>FNZ8b\NA0A(5,V[)A6acYZL59,[MTY8&+afg28<_PAA71.#Q,GD//
<dQV9^R[f(.?8e)fR>SM2(\XBI,=Z-Add#H^=#,Z]W79c&46gEB6=/_(W\4dMUPd
JV3cb2PPXK<Pe[4NbNab#LS(8B0WFZOL/D6/5C7U5N_Ub0R@1-P=]=8P@;V68fJF
eP2S2ZQ[:gSFJ85DLaY&6B,DQBLc92F4EPATGPaUH7JCC=L)2a0cBRCK0/C:7L^S
&I]E7-?A8S5LK3?cNKN4@&#b:RI[0#8&N)[CdCG9[-HaAObd]PaDbFOCA/N(O0,)
O:bJA&R1]NdUIG0cc?@>G,[:16RG<7)P/]V(Ea^4^T<WMR(B/UKF=8N9QF)BM[cA
ZU]c75-:5X#-6P9GFFYD?9-\R&+bLP[:98L/1M8TU?d0<;B57B^d:^eNHP#6QK.7
a@3)1#c?-fVQ)+JD-f::-LG#:P57a-5bBR/:F1CW^PYUT@CW[KYU8QRU-2EW_OLH
,&c+.N:aZC[1T\]J@2=]2A8X5RYFG(DPdR30>JZfWFL>FS7-PK5MHBO85URHD++Z
[cW@,D9F<cXOJ\5[7^-8+=Ge2aP.IUPAW5GbKRFN4]:Yb;4];4+6eCR]+f:H<H-Q
:VW4eIF-O/9(T8;_Jcf\-AC1-#9O4gcg1#S)@<1EDC,5VZU,6M:3T@FOA1^O#-A,
N<P(,)I[-9;7cff/XX6d5[J)6c[+HQ(6AO)e_CWaAA?P2X:]HRGLW]=-1(MRaLD<
(7</R^]VB89X7KQRAb^5A::?[KP>[3@1Y9Nf,<;MScD0;@c2K\6GK+[OY^?bLNJ8
82:RW/Z@[?HXRa746?>#UA=]R(,.cg1RYH)XUBUU9^;fLHE:bc1PMUBMW830R4EG
)0Y2)@KYMB6:)OWU\UPT1A=?7EF\Ve^0/J?143@B?)I#;I:#]^U)2&(g[HU[R5VP
,]6MP1d&c&F4,Ob?Ob(\6&N:8HP-aa1AI12@XT50c,:T6c2QDbSLIU4c\54SM?ec
bIB-FCY1_:N<=X\PY=)[0HYSB3HLZ8J2(4J#S7c2[e[Ldc8N<ZM,-PH)JB/acd:L
b5JGNNE@)0c1.B#I1R>dB3W8S>#-M#T<QEAQd06)<:8>W2B(1Z^FM\.ZO[.,/MPe
\fA,;3e1\eTYe30RG_DOLCcN1A#2C9F:af3QCC]0?C<,D:a1\gWN<D6[MA@>e798
JeH5^:)H<IE/<L&a9<IJ4?VX-:#g>9U2#?fgd)20)29M&1KDVHVWNI.M59I@4D)?
[g3^IWB8fKPLPMGV5O]HBdX;T)#>>?KA-e:fRR]BfQ?A+C;YG\VNbdVg6FA,-]IA
QDG^UJLe6AV?RJbS6A9:(Y8PM23SL89/SJRED7(=>+L#1FY/c@AR-E#E5Z=Q&6]Y
#22OIXEgB[TGbRTT\>M9XPe9DYb?I]f=H^E4QbcdR6IPAM1YQce>OG>7JP3:CF5R
DK^OS:aS0c[KB(J,H,dRb\?CSY/-5_cb_[<T>eQ7WN1PXd7/\:F3AE,PTfT)ZeV2
CDP4QJ#CeJ^EAS?6Q:[+5-K/:)CD]),&1L=[HNLI-5bA7HI21-c2L;<6eb[A(1TX
,IGB?(0c6_3+c.@cH.g&^)Y]d8,BGA5IR\GS/2AJMT@</Z3SQ)-#CS,:+eecd.>>
UbS^>B:3=b@Q;&_-F4=?QT89)13Lb@>&/a=WHKVb^,AFg[Mf1IOAfbRA4.QF7bgY
WCLYW9K,fL<-Sb;/DDgg4Y[;[d12fI[5+A+H/B=[@b55/6ebR##]0=GIbHYDV[ED
/5E)Af\&MY]Kd^LH1::>P[ZXa,7-FX94QIa?VI-?fb2.WTfXM<@)#,K1e\:(^^Td
F(<K?A&)LgET,J?B_K3:MWT=gJH5<XRc^WIV>38WB:e0Ub?X\>.c2bZ1V0P0)g<M
@?46=dDNWGUI2)@E)7e>eJ+@=AM=1S@1XE?dA,d+XAf]Xb=2(X,Z+=0F/4K>-.N9
Q-^QR07Q<AIPF,b(&64#3eE8_OGTHHbg/PWf2P<g\b-_5e@BNF#XC/P5Q6@9_\Q9
_V)c_]C2>C10B^^V3P&AI-\409C<V^C)7(6YJMZDTNMB0B),Nf4_Ad.8?M>.F7GQ
Qc.WU2I+AfT/<0K75b-;3bb;95^?>7/Xa_>19B\49]_Zc,3>b[G\ACfRUEc:c:d2
,TMb99MUCOeTXRG/=Dc-(-#I<:/92DJTL84#Wd[0)a-TU7V+(KTW78G,3D+VZP--
.:E:Ag84)MbB)X5)2J\.(V\ebSfDXc(GYK1@0?)6-QJ40)PJAbB@4M2VE>Z2T6,c
Tab/Q6#f)e9a73fY./1.cHZVG&+U2LC=A5I(E\Xc=dRY+-XC0U(N6I&(/2dS_L>&
1L/CP[Vg5YZdT)f29HAWcEE.T8d,6=GH.@,.O1BI0XNQC)[-(BdY1XOW[C/&@b=g
_NQZE)L3M:SdVSD6WfTbdW:#A5,JU:K9YZ::WI/KO.1Q,H]X=/[g<2+YDUS/334Q
-Ce<XbgAb^NJc-<V[JYR]6>dI:Tc_4/:^\#;cV[P@?E;cE^-89)Ffb[U/X8BZW+4
1.,>?LRK3JdB_797-FgH,:&;(D=,P5cQdIX3@1<#)Q5cf3^/HD^ZC712fRVUc;bN
FH0Y[M8K+H4((8eHGV/WCC[I]8F(R^;L&2Yg=K)YWUBgD43T4E^Z+a,JE??Z/72N
dLLYSZeWBPV_DBXfH2;S4Y,T71W&1:20WR(75bIC8bc29W9=4Mf6HFW)0EK=L)-J
U#Z@#d,_Ae_CbP?KTf3/_XfcI6D+@(9\U)V;]QU=3&E&QKd4WMaU-a;:YBa)dRI@
bQNJ59XBH\JA1NSJ0<R^,VM)10RCWc.-\&IYSC[J,f,O<O<W9)]&PMNKfOb=J+,)
?bB32?V^+@U&CCHaRYI;8P\0eLZbL#5Of71OJK(GMWgM.V)4/>a4RTVf-gG4JM:3
@K]1@2,407;<aGZ_IXZ9-G\U)FY?>X22)^_@F91>8_^+^9C(G+^YP,5+c-e>>[+G
>L:R/bBX,HE59Uc1#_NF[b9,2C^IQ+D[Y1Y\8VS@FIa.W7&be>\gT)eJ.Ig]UL]-
<MGIOHaKD.N+Z^R7L4\A0AB9\M^\EO94F9^:EZ92OD,&ST;bCNSE)Lc=S&KV?]c.
[IP:2GFZ=cDUdR<+44fECf#<d\c/g.2O(/;eWe&X;]4N)g]V42c7P29PU61\LS)H
7KUaWG\K(.De34X^@fL+T)SV^FAL_<M)[I09=@R@-8/K9JeO9FB,9\^Se,=]1B2A
A,QLVM360@&-)FVT.b&9[8X)(7F(A<._Q4)I0MB-e7Rb<(&S_@61-BPc(cH^B2G]
f,aF/^95UHX3>d:.\E,Z]?;dcV>J0C5-P-XH7;7PJJ64M8cXR:TYO7[=YPSO0H9S
F]K+P^UD+ME0J9JdF7S@4?P\W+KP/SSWg7[;3]ONA)M^@ASES)@5d_HA>Yb;.Q<,
;?X[J]4R8CMTfTYdD22=T@3[A1dA#<0cO=@3]BJ<L5DCeYK;YJ/1J+c8B(b2g4OV
AF3V]Y0LB4_Qd>8J0H9D4&Vc#6\N@IRBJ3A/5>&HH?cY\SF+,>MU^OQfBJG25&2+
&g4g(M2F<(fEE:P_T^g1E]I;SZ:#0OL89\:MT.MA(P\W5<=OG,PGAf#_-74>e[UX
+3K<BQND?=6CG,+1CMTIgE_C52-fAH[T^/YIFCA<g5E5FgH6@F)Z-#a+^;86)\d9
HU9^H=Y6GAJd6Q42cBH>S^Y#J?Kf>KKT8f0ZH9BF\\>@[[dOeO4RRa(Z>\W?9?O<
3+TDb/]<\_1-I_H3-3,BMIXJ+gK)bUEO<=G/beFKD0IF@-))PaRHaBE8)6#f[IR>
XC2bOa9E<YQDfYS3TIK0W\D(?<TF+UJg5;23g>b]R04APAdR\ZgVSeL;#J.D8M+]
=^4X;T51N>C@9?V)D/EQ54C&\Uagf#c^AS\O(/+7#/C[@84+2\TTF_WSGAAFcU):
dGPa]]^,DB=b(:\E2MYNY@8Va+Q-/]_F)D[I,KLT-+VQ)&CcE8TE:EUaU49,dAgR
SBKFS(,9,FC2;MJc=W\<g/PRF9<HA3bTg<4dCRU=G1\ZAO<9DA\&M<I;>GCAVb#K
C1OS1VC]?6E9?M/cY6(,/>4Q3/S,0A7R=B3+4,@@cSBS)<S+^f?cfY=VA^[T@eW&
\H/#f^Z6-gDECA[.,_F0CNLEH)7(SHE1OSW2,=(1CPGP?)5K<37Z)&G=+:>8XeE<
9QV2OcM_Hf,Ic@+)C^bJ<>SV->9PF3#MG613SP:CF9dP\cO5#dP8OFV0HMLF+D#T
+fg1e\DEH5^[C2gT]A[H#HPJ6d0-1/UU_,-I2FDEEF.,9>)Z:ADOZ-M;e<^c8H)Y
?2Z>+X[_M1Q9>&1bYXI=+QQ)M>AO,A8UK1ad<H1?A5BR(VRD.@g&PN9VTA^be.J5
KIIP68ZB_H<@\L^D(2&8U_9ag#>UJUO;g9A4^+a](K-JU=O/C0#.F1IbDEH)(.\M
[c,5gd^SVIbIV2eD&6X>J6+c[7&DWW9Wa+#<8K@8[)R:E2/dD3.ag+D/ZK3YW-B3
1V\6a@QYM[H-YR1>67-eaJ0f.Q6T]>Se.FM8g[E)=>WG+6cZg@M)O:(98J=#1B8^
.<43Z-@36[O0)KcbCFE;A:]JG4ATaa<f,ZO5;(>Ia=g7S>,2W0&CGQ9A#;a=CK8+
)dFM)8I,bM51.Q^g+d11HPHRUeQ4B(B0S2BTAcAUGaY28I5Ve3aTDa>#M2@>Y<G8
MbUf[[bL=)>_>V]+K89MPHgeEX57UPYDC97:Q\>f\gL/cefKXEZQ._.ZbHPJQU-U
)X9WD/Va5GBWY37WPU;LU/JY&gWdLX/J4fW&==U4A5cO@Ib]M:G;JOI[98NCO-.f
T#:,[9;0UI(_HGEOI2#<PT2Ba#IZ:]b<_b?/WV9ONV2^7;VFN(:JJEc>K<IAG1+T
HUc@@a<R],@/Z&-0:ZF:1SMZGf,aNUPHW?3L>)fC>(_7W.[=HZQL<Y=YE-?/Jd5.
)RCDCA00Z-<[4[F#[-C8EI93L78e6VDZK@23@X5BeX.S#D2LHRNZ4;QdKFYdSge&
N-LgaY#HC/PGQK@[1N&B?^SUHVMLdT\6@PQQK\3S/-4SZXYRL<<ZS8D1TNe_O6XZ
TBB&YWG)/X/dX_XN_^#]O),c9LC>FY9F>da;TRY^Qg<-HP>Q\V+993Cfe^<R.af4
1)+CNI/XOA?:Ga4b_=W]O+\ef);)NP>KdFBW,IN>MCc;gVHK123e.U;:>W?ZeF2O
aFa:I?#ZUIU3(QE\4.Ne2&CaZ>APg#<fe2bL25G,3KAQ@#2H.;0;W8WGRB;W4>=^
7f/FLY#<MOeU)<^)U]^de]-/3CXc.fQUFXVC5CX=D/#?dKWN(#Ld&:X2dScNHIX7
GLb3^=\?#&PP;UQXO9CN(/)3d8VT6aW9?SIcXL[B_#H?[G047S[VE?&M2J#=H-P3
S8B,,e_1CYQMa,<7IV/&.2>M+FK==(L>NRQGU.#CW[CDC]aeTI+YI1,,0KVTYUS.
+Y;B=F@f(Ce:.gEgK_96B=T?_5X?&,H?17]Z/6)F?Wd@(dZ+b+RAC]K;a1]P=V&T
^b)Ld):;0cYD[TfM>?SOQW&_O-ISW;>3)&JDN\a5?4SN)H5?5BQS@+91<)L4K7g8
#CB+-6MVPdR2P+I4T+T6RERFY^U9FML7ba4a-4,bRZ^[:Ff&=QC5^:E4T\)-M:MG
I,e&N]dNOD2\SfP-^RP-e0OMaB:MXI@41])><]A<cXB-Q+<K=<:;+?fTbDEB.K/4
0:-M1CWMed[[)Q2=cC2KaYQBZM1X=85YGVHK:N(5A-I)]CES_cGN<AN]U2Sa3bbc
a@edD4/OM-.9.013KIJLU3\Z+ac5b/#(2<.;=9H\XQ+XQG5FDE(=N4FZW622IVYK
(OZEDB:<Qc+>#gdg/f6PSU7\::LU6V-(</\.S\I=S.QRNGVB)PfH[9=,+E)#-g)0
.)UJUH/^9bD4J?90f)<VX-[bV3F\JP1ZQLXLHT0+<a,TSb^[J,TIB]IELCSCWX(T
^P3a;PWWf>3TQ1Yf@aG[V;EY(fK50bf9XCDKF.4:#3FTIR09fF8G7bXJQ0\I,T]S
#FDgTU?+K,XUK;<V&2PJF=>R<1F#(IUVHPee0UU4^+R12CK?FCD,]EGRQML)Ad25
I2YL[f,aS+?9e4T3T9IQ<g1\5Q^DG:H,Q7HAJ:OTeb<5B)c?HNdPf__A7gTfK>46
H^7)RA&CE/De,PE)XN:dP?@8LA/)U:[e0W3\[.[(5Ve1F&XD/>07d)f/N]?&:OGM
0CP2ggUVU&e#A1W@/-:RbW,(^)+c9f975>3\=WCF.XD^JFc@MIU-9C7:BTF=W.^2
97Q;)PVNQ[Da]5X1Pa=Y4C6+_4MX[3WI5Ae-IP4gWX\G621ZB-@NFf+O>M<8d-R]
HY(R)8L(W<4VD?7N.+IHY6@?\J#\eH&@V1U.WJ()14Q48^d2)<gdHIG62V5<G1CW
DJ2KE)c(LdWAUB2aA0/+3P:WTMX5-N;.\/XPQg&R=Ge<)Z5MgF+ZDV+(4T.[&c[8
-cZR_PMB4+)YbHJ:-a<EN6GfHQ&T2g<D^]/MTTRJZCeSBI3gcf)B44Y+V/_]KL(H
#9TG66f[IRS9-=_\_Y@[K]&G/aJVECL1N-\>X=Y_),>MC;?W6@5J8e.S2bDeXdUb
dY2L4XVLeEc96P9-@OJUMET3TH(U\ee(]7aa4?K2?I^7;K;VaXK9OHWYLN?bg0[e
OC+#+CT)3>,,W13</6KSW-[4df]7g_SP4&X/0SB_dK9/0L-#(5eANb05I7RDRGJQ
UFS:^Od?@=L&-^g0QA&-8O-62A9\Xa3^<7#ZVO2/a>Naf\\Bg0<]aC?NIEggg#IU
B]APDa1#5:,=0_=&I303L>a:Rc;P@\JSgO/,UQ846VX.BP>7@+Hd;g]-f3.;U7NK
3c^V_,/QV^U8@[LEJHE(A\LW.].+(U7&E)K76MM:95^B;J(F=6\L.4=a\GV[(NGQ
WNAFR^LP)YN-V.[@=WB?QO8Xf[QEK:HS/-/J4F<C1V-f+IK=KL2E)-^@-5B<g#Z4
TXG.Dd+9NF;>E]eF\C[O7bC\D:F:_:T8ea4&1\J29JCT3SfbQ&^^E#Z0,7+3>?D^
&8K23+-Bg3@>HdC.1V2RA87DTBJg^cQbNG:>]gI2d>P5GIgQe/Q1W\Od3^9^G#,Y
[-Td]@C>3d<.c0>0R8^,KRCN:>?(C,:9?\Ba>]+0cP#8MHQ[3O_HV-/9IbVMZ2eS
<SZ_>1Z]KL,5\F&+D98Bea&TH@JPRFVF25ST@4ET>)EDH?7JJ40Z>;0NIe8>@G)3
A>Ig@WbdL53E.;UIX_42He8ZX65I,<M(3<VMLBaf?NMff&W?LYVQ&ZK+.e4#\WU+
Z_PZ?IY/Za11KMaX.?T>=^]V8Q<S)/:c:g5<ccUD)X4HP,G.2D+,;Ae8:1P]3:M/
gf<^WO-c<P_Ze0_U3IS^)R)-/EY8._1d76_LcP+A,Z,B+]dE9_+E9;IYL1.?1bG>
_@J0^@?N9>&4>>OC:0OQ8W\&/c(N_\6NdYgI0X-Lc#YGg1--7HM&eY(P8V)&U/LY
1@3&f?#Yc?R7SF0aDKWZ0[Pa,d_,@L2b64\/b@7gWDZ+)(0G9F>BR:J8\NU-1IQR
?/gP)](5F\:B23]VG,)3aBR)aF\BU?c:C3>PF_gB8L>7LP2gGcR?X_5S-B0gg:Ce
9J\SFE<>MCN?]=>63/gU?5,?/:FNJ,;YZQ/g7[26>P@M<CK_O+YOHQ3^CIZ84-YT
?VDd+[P(e//796RK?_>aaQ=K/>C69TA?1W8V(8-BPG,B0eY[=0Z2B@_81P+N44Z:
CNcGKXKPXM&OMd8.]X#?U4)(d[a<UR7TF9O)75;Lb3YCQ#.B&@eG+G9?&YVg\&DL
>Z/f81I.B_ZO-EG:=\R]XYQJB0(BD&I[>dc@J-5gb.E,^A_TG)BV0=&(a7T,]7-O
=2a<X&7adB7_?WV#IQY<MV_^Y@RB-Z/+;1&=-/>G\-N,=-#bWee[,,^ZPLDa1b#T
5cS(6:CGW>&GC]_d?=]9a+f.^g?3Y0G818_eY.258CTX7#YdYQ[E3Q,AHD<FA7e<
_cb/J0Y0f^1#3HL.@I.fPF8c?_ER[GB/:bE\UF)N\Q67&B,H<QVQ4fM=&8g#KQRC
6Pd6GUe&R;3]8BXcc8?([;9?JV1[H,EVf(Z;T3A-D+D^6:?2#gdL3;^@C4+VBA?P
N&YH\_eJc?W@]K-\PcgDTe-/E\-dC/,Y&>AK>?;);NSJ5RaYJ9+ME;ZKGNa8JeEN
]71A?1Y@\VUAM^EX#YeH._3P.80PF&I02^SCXc8G8YQ_Fag[+8LP_?[.L5g=><K^
57ZM]##T@]aME.HO_[QR0&Q>@f92&:^S41U/;PTNJe+H/C_>:+4GH=P9c8?Ce-QN
>;d/&d_\9=P\9XE^TbB><;b;<6Z^dZ35;<.adFK7[WF+-Xg?8^,3L[/g(1Z(FU0D
.\<XN-@WXfdb(ZELc:?#8[YI)N/KX317gJBWdRQ[XMaB]b-T8\RR][3dWR_0;ZZ:
Z>Y1K3;,&+SaMW=aeNf;TRR?VBYH^08IP]Q8C#6.-C/@#JU)?2TK0]-PH,I/]X/Q
f,F@Wc#Z^O;\.N\I4)&<f2[1^CP_^3PfJ[-6+S2+ZCT#JMFS#:OO)MQ?TBWM^GBL
XV8<PUXT>T2ZWc@A&GM<1506d3^M#PKD]c>F^.aV,-]\4A80cdNK\14;=-#&aMDI
LN?_-[>T@T6ZDg^R8;0G\8(=Y=NBf;?9)=&(Y@.R-@Qd41I&C8PR(SVAIYC@IZ+S
a7EB@F:2(\X]V^73<Z2LQJ8DefaDeT=6?,<7b0H8BL_)Q+6QJ)#AVP2\4]K&]1K4
>8DB:gAZ&Q]\[;7)-93G4eTZ7UF);]_=V^KV<=\F;?/1NHT0;f6K,NYT>X&7MCMF
ca]CNR^FE0JR_#<3K-4W8?R7N.,]^743;1<0A?fEWSRaYA7gP5L;EXbB=0J&6()d
27;1_QHGBb<JA5D6X\UbNVGZU),071Y9>INN]bAKI[O&)-,]L-&+G/S<g[]?gH_K
GE]XBd9_-F<^[.9\]eKMKJS2?FY77TT5NY8E-2INP-Q#cP_QJL8-7U69bZIZAfZL
cIKQAP:;)UbQ/-[O(HPEUH4W#/F1BYZE<7I4WR+d&P<3MZ<2fT2U@@gQ:=F1:,>W
Z_8a?]@gE1@KfN-].OU](_1+(W[63(Ta)2TJF^A[+e)e^_D/PEQFB7W2=aOEQ\]:
>KIH2R_>,NM._7PMg)RZZ@4c46KM8:+b?fDc#X\?dEJ+0T6:5A)a-EO@.A+2=<8^
X;]G@;2NI(EM^VYG8J#gX>=VMEEgD8#6AX?S9>;eM5MQX=@+-1CH=G]M.9#gB4DR
QV.1S@K[&PE9@9IC1X9_2LLReUX17[1(EQLM57ZM5=+8&(:5&1_;CCC-FPd\MDZD
B01>f&^X]FB\]1CX_,Q8@4KHXgg_8\Oc(-;ZBYOZVZPMR0<ZAA5:WM8[C5geKJHB
D4UE@=LDF8]4N[=[E<d.2<a?I>,PE3[CL]:-59Qd=-[EY527XF>:R8&_N2@OCGK8
#6DJ.12G=/U-BMS8GORE1PJ/DML0^HWQ0&@/TXH&ZJ569Nae5GN7GO+(Z94.,eBT
__^U\Ma9-:ZbIfZ:..P6?6RZ(79U@N02bZdIL:Lc^gX#P7,-=2-(,Ug/@7D^e:gH
e]2K&BB747Zd5Z1J23a)F/Y4&F+[XG/DBIO_1?2cgA)6+@V<RegM<g;QT8T2bM0g
\g+<AdJ3N@\;A;/N)I0/5D56KN8Y8/<c+Z74Xd93b3P3aS92@61I&C8Jg1GfGSYL
cVA/)7K5:)MIG9T^81#5.L<bP2E1,62FA)cTZV\I/TOfMU/M6Uc]IfR(1P1P<#;F
\NCI/c&)=TP/:^MU/V7C^>)3=[J-<(MB.&eO+gS5:f9_W.Y)>KI,C;QBR4=FV8/Q
gYU0Tg2g_RHA/.Q8NBOUTGcCScfAfMKSPB2Z<^5?BFRN[V)X^gI\.08M6M?HCX-A
a30,BES0D:,=Y9[N<Z]UgP:@3fBXZSO1Va5Y(C0f&Ubc52eHZWHX8A2a0&)&E.8?
LMA.QUd(<@(7_WB1@E+<-M\g#dW-^>&9T<g;JPQDT9.c#S=_<I^78VJ>Yd>ge5WY
GF2@6U_ZOJSV0[M22]WU-B8-]#M28[MEKDT(\fd38N;?:O95&O.Z4BbU]9/EaJgF
YQG)O=TVRLU[FfSK\BS@)&+f049Bd<d)CdABW6SA7Z[Ba=,DC?0?Z8)HbC=.8RIL
ID?3N_O?BA:-VKHPYYV?)SgJ:WgNI)I:,)N.>-W>.YQ1J^7L\E2SVV.Y@YD__Nb@
A3Z9/f<<S92.0;KSN&HRJ><LKT0d];AP\1NJbB4MUaa\&E]9&6gV7L;9fJB.[080
Q.WSX3;+#^2QcR3e6,Pg,>+XR7Yd(J6+Y07E1IW(DWEc3BQ35@b>ZDYSY1/MVRO=
.VM8.>GBP3/HG14fHD)^-ZJ+\J36<FWfXe?e5SMT7g[fZ9?\(JMgEK&D7C^F^6e(
>SA]ARcIN\AULcR)NI+\=#P(d8PLVW.B<Y;>E7;Y:F-cG3.RD7D/]=X1O0ZE1&SP
Z.>]dW3AC>GS8=3:Ab]5/N))KQFf,FVHAe+dB3N;B&Ve2?E#6\@#.90f<KRfZZHW
aZ;:cEbefUcF0@935J[+-@O\?91O28(0a^+4B1/e=GX13+EA37]#1FF,cM;L)+PA
d?05d[/f#E\+:QJ35Me@)\,H&/T^H(g:+&+X8gT?#+UNE]bI.DfR4<ED.[ZOJ09I
Nc=4OMML])34(:Q<>-=Y.4f_&J@O_T>[f#,GP3-LWf:cWXZXQ(@IZ>QY?aZH:=2V
7IL6(;#+BV0)Y9SJfJI9#W:7F[+e7#N^_CT\Z)7Q@6MGF+Fb/e)5VC1cYY2?M]#B
&FJJR[S>?TV^g&KZ,4=WC\OWT0/\fS\^?f\8=C&ge)(C[QZ@+@9Te<Y->-3EaRJY
U1EXCQX@-3PHec<>2]Ie(#]ZCa@C=5@VJ\W\9FTK^V]gWfU-LT++8Q.VfD\42D6L
P5(6f#\<SBa)S8)GT3ZR(12<<V5O](]LHT<UUH70(.1Df?^_OG^P]ceRZ5<A+?&X
AAfR478VNOf[A?SfO8eVY)?DX[1GK/VT.0CXL-?f.P+?B&^W]b1-IC_KeA3_-CJ6
+S3-3_YWN?[07Og44\-b90e)M=LP^T>7NRF4;CCdMV@=8-&@)VL@P7&LS>U6&G5E
OIW8O/+(1e^>=&\/g<9;_=A51-F&V6:,=HT#gO4^c&MS(:cO9-+L@I&P>P;VG0=(
B/0NRFfeP7bWeK][YCN+bGI@#,3&@+]44=NJ>A3P[G36f&A2.+2H;(^,2=O-N3;]
.V^0]0^K-T).P2)B(MR9-HAT&N7QI)@FR>(>D3S]_P6FaeQ#VTCD].SD5#.JgE,0
HQa9?B_<F#S]31b-.,5]RZ/HBN,5N31DdM?UR^DVF[&;RRD=5Q:D66g#cQ+NL]&Z
)VJJf]M3&[WdGH.aNAc)7e&-6&OFd2D+6][Mf:[Qd,WER9UAJ;Ge7cM5b\WS4H&I
,2BbBf(f\G,2-?0U/c+V++>TGZLK\Y@CS2=P;I]B27S:=FP.E.a31+#gI5S?D-?I
C8QF:=D.Rb\>D3#c:gF;;(]Igc=I>cP=OTGDWdIAGFae,Q)\JM,_O/U92a0f-JG9
.#<QT([BKWKOHO[0YEgEV,3fO5T]c-U-N3/bL7J3R,;dUF3ZYTC:8N.NV8[d-?Wc
8)9DL](bSMAV-NUO(:9FTP[OXca?:0dO5ENW)/3SDQ5Wb,ea<.cUBH[@1=D6Obgd
g-a)R9O;S[RGeBSIa4IWMZg]R0,VaP_1-.:-G_4XeE/dJG[A2KP?cRW<Rb^?YR7@
JcbX^[+J?580C3__/1L\K.1JZ-M(_J:TQg&.)61dV0aFX\1Vg&KY_aPg6cG[bIIg
Q@+Y6^Ce+(9-6,SPR)c7B5K6YO:U:1Q_^KC-RL_A,&YT-ZZ/OVUTdU1a:70)WKb[
AB+GJ2Q<d>L,-1FYKWZ@1Uc5N7N04af5RFY0BK5B8B()P3dN4](#_dJRL:Wc=61X
NNGU^LT+@383S;acbN\:J74I4L=TLLM?IM_Y710Z/K0+I(0S(2_C#TXIE&@J9J?2
?Y4HaR+1+4@G8&2Y(J^_QEcOEegY:3:(&Ub/RM<)UdabEGV)/\47;(IX5V0Cd_K2
;XPb^M41RV^a78Q3@#U;YbUE2KO10@HYM#,:&Z#1R)/GL.?Jedg5AdR4:fI&A6W#
KM2CfP\X/<]RQ#eXK6K-)dUX+2C@V.48PY;AQ(f,]]KL>H0dQM=DEcWU0_4JeQZK
E;KQ<(a1H;8C80PS,F;]^<(,J>I[gPO]/9@\bK?\/M,<02g,P@)aVd7F[0MVS/+c
Z#99ba,01]-#BU7KT2\-#X#IYTEc=Y9C]c7FP46Dd2\(\SgeWD4<3G-SAJB]Ce2U
#W3):G]OFJA/f5&.8Ig>UKZV2d6/<O9&g>)V@0K&^S4D]6(+T)_,S+)^1K2FM))&
H[E1[KK.0:99B#\T1fJYNBVSC?:;8>_4a.?\5KC53L@.B=Z]fd\ATS09).>13)<a
UX4;XQdSR[@IIdEeON-cP7C(9</TN+d_Y.HSX7>Q#(?gB[K>&FB0[AU5ccKIA9_@
=Yfdbb0b(TOH6<&gI93DYYRFS^7e9D,D-4Ab95f7E@^38Da\E:B=@<\9GeF@&,U?
XDS.NJ2XT//MNH/IIA/a\_LG@@XJ6J?g=AIT<I=KM?J.OU.ABO;ZB#1=d>_>JUCM
_d@7@L?X4PS&f;.(KHF2P(::a:fX0fPGZ\&K1P@]fWCZ=CaLUdg5G@ZdVcdaU\B\
C0\=BF,-I\([=bW2UJ^Y(#,>]<[,cNFC4B=;SL[W:#B.1fS0/A?(+_U5+1@R/:&W
ACGHBF&Ne0f1>e]54TB,=7<?GcG+g&f)NB]\,^1aIc[9fL7?(8@&DV21/=f#5QN/
(eEdYc@=[00.^&aRE+(QU7)BCSgT[^A7&GSeCfgcZNecCQA>MMCbf5FQ&EQ:8Ze4
cbd?N5fT5<6+MP]-)Z89G\G#=Y:T\H2,^[?31S)J(f\dgAcPKBCX>cDDRT0cXVE.
CP=ZFU6R77B6WB-I#<ee8L1@=NJ&2@<@V=f]?c3a;2R394@2KL:eaLa09=eR4([?
K79HE.=.]MV&8U-U1^D?W^/W(L1R<aZ9^R2HIbLdbTT(::\K&a66aON0\cQ3<\DK
fge2JZ>8MU[LBeV23+a\\#aJR=Z:P3<J()f=K]3F\H[&S:;_(<VF)8C4B)OZ3-J^
,5C@5,)&;^K,W/KT&(5M\FNX,_N-77C&XgE#Q4AeTUB7XCIE/:4cUL03]O].<8E@
=GS]&5VbZb3MdfN+ff5>.2Xd8<81FK2US)WL]YP>AZNE43V3d=)ES]D0dGQgE]R_
<e[FL8LdPG_^[G[//FBS_-MK1g_4QLRMT8OXSCS[VWf\[]Mb&WZLJ9<YOf:FbQLM
J;DKR,Y/77gBXTcZXTL)5=N3>7e;dDH6J[_H0>)Q_53YIgY65+PKRN..)D>;W_Y=
3bOSJ,;JDZ<ULAA2#\D/(/KE+M@d@DLYe/?[C/[RKMf2?E-C@I75gO?</gVC..3g
Q(0GeaWXM9I;S;#ADORXQ67dd_,Q?cIgO2FY6E76/f>B7;-823??FR:WQ7]RMAKX
0&>a>>Md^,+OOJ^IEVXK]MfJ&9837[Qg+INEFbVP\5J0dU4G7][O<94D4M1bJ<bZ
ITIMVY/(DfA3EK\GAJcQM9(:Eb)f3R1LXGK@J<]>1QHG+,bDEIF.T^@PN;NU+[4Y
V@abeXXUT]bSDcJ=RC[T.3DA&.9E_)DPO<(Z(eW^)b?FO;ET&TD-24_+Y7A&^T(f
,O4AEBeESb1I\X4b1WPJ362BS^?_b30.bBGfH>deVGHf12G6HPJ5D=Rc]&@-BRL3
BS@c_>FA)AG]K\:MQG_LV0ZO9TVVTTX^DM>3\B78B4Q2A7NW(:c^4&Q;J_K/(&eH
L&X8[;CXG^N>S3=)LWXY=)_@-b.d#[dBBR4U2JZ^L37YML0KEK<<R]f/Ge[67-OI
fA.bUDX=B(aHDR2V2\K,b,G^9>OBP()2:>,eE(,1Z1/^PJ3YY#/,NG@KMO+^QPR[
^-KXS8#)Q9.P-;/B@fJ>5;2@]2J5;;H-8TL9#1aRZUZ-AdW8+?Zfa5]9<B&_ed#f
<3<&E8]D+A]NLZ#SATA.V#D]c^BAK:B2@R#^9+IOPUYAYD\4-#c[Z)cBH93(SBO@
^K)39V2L/DPH,G\HHbZ(FI681Ae1&\NN+O=1X7K:X[JU(\gfJB:END3[O&ZHG-5S
_Vg>3DfZ_WfFaR;@E?/a4=L&0QUYLU,PDA8X5I1B[De5LV9).O08=#HCA=:7d#HT
c=OcW+6:f]6[-/N9P@Q+&Ob&5Oc7b(H75<HSeZY.b/<?;L0P7c9XHLR-3-YY>SZ8
H>\VU[ZeZMeVR.3QBfYV:3O2)V.9///2)+\YQ87FKXH(,AK[S2N]f?JQCOR1KV,#
,V[<cH_)R22PGAD_WZ_?^;DaF7KT[5H0fTV9QeOVA:Jd\V(WM(#eZ2R8++7^/]0W
0GIG1F=M,dVFABcDc).88RLCfMf;VCZMVe.R15>,6O-=;(EA>3B@T\eVY&@7g=c?
\(g+F&N<=bQWE[8HQ1@QTg56B8F(-A:6=P506)F.8:M_)5._T?S#]T.7.cBcfO3I
]2J81KB^F&JSH.K+A&MaP.\,G<SK8-4:=\I&TG>Tb)<X:T].J=2gEG1_^;dSDL\a
\3J3K,#C2AO[CLKZ>^TK51@dUD1/a>Bf<FGZK]OJF]Xa&7@OD/<R/IB)0;XXUCCg
Dc6X6ORN.54T_EVP&Ug04TE:&3;e2K7GDAP+]07C>Le42A9_dGB.eQVaI[JC[NME
6Q5)9\E\KWb&3;,_,B(^XRC^9_+1?;L+?DNY;_26+O:R3@+XG^[_9.BW-ECgLUKI
VB>ZOgI1E=+NO63@&/ZMAc0XbXA;YC36\><(X&,1Z5M0]#\TO^F67ENK(&3-ec+T
>QO>(-eV9A?3AC-e<eLWgg(aU^4[A]&OYVIS]06cJa=HVa>9\-=D?.2D\dPeUDL\
=83[.B8RfNW(7=DGB)AO,XObZB1PZ\Qe)B<8cV^.#&[)R[G-DNEJ7HU^^W,??SIU
UI:FRLeL_9N3E7Y7eSPHF2:3aZg)d;dGb5Og&X-T8>VOKY4<Q(=S[d+U(JOKEe+V
_g49&7&9@G<6,U?26gV/#6HGgAZ70WHMYg;=.AM<EQ(:X=&4UNUNZEPT1_,Y8<H/
([G4[#,2>2NOJ[:@BU?gPH.GG+cFX[#L)2bLe#B8f,+O/deP>6N)3H(:&B=HX@Z7
5QAT&P)5M)/=05#+Ke6fC:D^e2YcHW&BB91X^a+Beb&G]OP<S[8EXe/F280N>6[g
_K5WD9]U7Nf>22UNUL&G;;4YF1V-3;E[/LWEMT<@#+6Y1;6(G,.WcPH_-[ARO;JS
/dI\H4,:gBcD3c0#eg,@[+RALS,WO(_\BB)H2A5B2RCK<5fG#^M[-68\PTX9KGDJ
-1e7.Q<5(Ed]?N^S4[WP,)X,1)SI,g_D?NLbJ6H8)5F-fH#OWOOW(3Z(Z?);,6J3
L&4>bT29-#C3?KKC9[JL;SX]FA[BHR588_O^;D8P\KaEd-dXbH85ZTSV>==+Z+IK
JI6KX0RbCLD7H>[L,4\IaE0,XYH(]SFZ=Uc.eT(e=2c<UTY>02-@U5R=@:0]6gWF
]<T+<@bPdEI1Sb)bI<[ODM0IBfDMN^NB\]ZB([134([5#OCdCc@MDg[FSYU_,J0M
V=4L;J7/[OW/71-_D,/>#JLWYTD@H(4YMQ;VWLg)6KcT5YJ#N[U0_c&4^8PL=2Df
:_IF8F?IB:74R?S7=MdcHJ&YK_1=[H&1^Z/TPHXXVQ05[f+HA#DQZ(.DW^YKd,55
W,VJ#T>XfR?-4BU>R\+,?e69]OgN[317ccD&?I+]__2d:OAEBQU+M?E[S84CeY<V
+O:GDM.0@cf5@E-?H&VXg2/B.,+4W]Q&LOFYTO#S,DM5#^egA_AcFQ87Z9QG&;UV
8a4[Kg-&^-K<_D2J]1-c6CJSdE(4O-a;@]>B3Q8&UJ8<PC=8Y3Y2.f:QgEBU\>a#
:d=&dfU^)W:VZPbPCS\gH998W+2FWW8N3W9WU8#/K90G(7_8RF:=M?)A88>M)5Y1
?RW5I=eFLZCEe]QEIQKe_fB9[.G1)XQg]T:C2.@]ee^]]#K&57[YYW#\WNY5gZ^b
4>Ce;>0ba+9,/^d>+EbM68PJY0e=1<XPC]]O<QV5QC[834&TV^&\HO1UcgFG32F5
U.IVb&T_X<YX4d9X4JYcgR&/EYG=\-4V?,-(C851d:]dXHe\@a#4K<Cc<,\eQVcB
\3FGEUP0g<JOWYW:#MDcfEMdGROg^(0H]92)<X^a(MSD8WI8b.Nf);dNaMIQg5?5
@LC;6CI+G+R3&BJ8B&B31ec)4c.fNd\GX8-,N07BgcS;AMXeT6>D57[O(H)^D]KQ
LZ<3W9DUaV)^<(?9;M=7F#c-a?/EL0E;X()d+WR#/99:M;:BOQe=U<>fW6I57/9J
I]BNa5HRGBB&7JeWK.U2GWYWDUDKAa3.2-U,<(5e,).Q(.#1VOZ43J1(LO@=bWR+
:=YAUW64L[.C;YRI4>VRX4N0_<+5PD&GR]^S?B/@&P+MI1Q@H7<<#F7@W@aT-^6[
MY1bOU07fOCOFKVW<aO@b8LebW5XB7/\^KX=#Sd/PQZOR-(6];JM&=0d5d6.04G_
g70>cQ=FD7DQQO+a>7+0\>eM=<E4Y)Z_MJ1f3CDR@=Cbg=8Y^9NKe]f0P53SDI>M
dJ#,/;f42UL4b,cU?KK\;Q6I\[UWfA)9+-(B[XPM&eUF.FgMKYa1^\.?GPB-4N?>
,fCV?S\@FeK87ZQQ1c/V50M/cSSO,aPO+6UB(?SZ-bPKQUUg3D:,&\H[3f)4(,&d
7b8BZa6::c-8Z=B5=H7G]WF-/[5YY,2>^/D->Rf+\8;\\NA57.D@RI+=-QY4&802
_P1<N8;IbA_=,E);[3T.]aNY8,EVa4._X[:f_LGHT)GKe)\=OF97YQegTG1&IR\#
8OIZ^6VADQ8(b<V]dVdC14A+,56/KVe<FOFB:N6A;ECZ<ET.WIVL:WFI8FCO<?ab
g&4VI)Mf)MdL\[D1-<\.J\/D.<SR)\O;O3FdcL(fL[EcW.9a7Eb]\Y4A39[+@VCB
Zc@3Z=+]82b8K4ZOda^>P/)Q_HO5-5.c1NK4F8cF8EgJ0_a9D0QdJcUg]N<ST\bB
=WLN)F]ELHXaDY5#gFLgP;Kd2WZ;ZfR<^gWOX>/SfZHW,a)DNQWSTKXQ9U)Y/fM8
-.a;dX6cM[P.M<AM^D9.5SWRZQP+FU;H??.d-?VeEC]3)ZN)MaKZY3.#ZWOH6U;b
(XH4O1Ee\UO]>U+T.PE80H)I#-,gC_b_3RK_E<E30:F&QI;FIZ[-3f]E>DP@&:?]
)V85YZ-S=[].<?X?#d6(1D86H=ER@+X#d]PK(RR91X&3.H/H9&-5YaTe9)R_a<@M
+6<1#dOH@(_P18SN:5O8J_JM)8@IQAU-BU6(16C#84&W9>gX.K[MdY=6O)4ZS;HJ
ML<?6PK&@Xe5-3UTQI5L.RMLU;&7c7<SX5:7@XF8P58BB^DZAS5O\WGR6<3[G_(>
C6)dQYZ13X[Z3B@aXPda(#c1;Ec?4)UB4K^P4N4ObP2G[M7b-d(cBIC3-c4_/;#T
S-Zb:.IAKPJ3X^00)Jd@WfP0U4Z1&^>WK-E5a;J;ZaP2B:<[ZOU5@\Kdd:7R1AD4
4Q]9#-ZXdAge=U94Q853G;/YU5X/D:)-2eR#>JRK<^e7c&7Qd\E0Qg@#fS8,e3+@
8OZOHA6F4&=D<fYebaN2M22E\9gV:2(3@7eEY]U&Y7AK60_&0Y[\6&:67)]P-8]S
,g4EGCXK1SB6(&#[LIO^MddL<W(NU:O;C(b)_RPQKQI?Ze[O@I=7W<49_#;dCQ.]
<BccFY:D+4CYM5I.aD..@e?acS(S0a_[8&Wg9O6POPK)Ng.X3HOWU>SU>R1K7IVe
g\RL.cS;_8#K&LH(KT/(>+\Fd3\].6Q-Z^+5^,M@.FOc]F5V1SU4?6:>@B1+G<Y>
<E^25+A5A3D]1_Ice(+WJ<b[8&WaQU_140<3=3:M@TQQPd2cPHE&1Fe[:<X\f#Y7
W#K]5C11:=K+e_eN?FT67:<;GdFR<P5MOLV66(:CIK5Ka@S3bHZT7Uc#1X2Z41H-
N344c7M)#;<=,NB]_\.eAb@&<J3C2L==(DC]^))g4_A&W=+)@9^B<@^RC(FLJ0BQ
gLWNTXS9\X8T7W3e=7UU4<fL.2KR=42FgCTA]AFFXfIL8Mdg4\YPP2fZ5WTOWBC9
9P>)dSJD@SZ+a7L>GZ.-^+XW5,F96+a<2c^f#/[,^b?SaS,5F,)R3f[NX6EVM-E=
:US<W]BV4(IFWTf-aB4T0CAU4.2)0YgV5f,P<W)aE^0c@,NB^E@-RET++8V6f,BD
#R\)K=dCd]@3DfBBafUK]FFe6b>^N2DP\g9SW[@dEaX-1#88+#/Y&3YS&YY\W,SI
)?;N-,URG+[c;@]GeAY(:>V#4(b(be-\VAL:?^50=K=KDC=CI>XQ0U]ReB,ZM;GY
9(dF5<:0ER)ZEX[c=J@)EX&SPCO?I30Fg/VL8TR1a@.R5c2IEJU<R0Q];B>PTdJ[
-7F>PXZXQ(c:N2+?.X#(@4CR\JbREWF+ET-O[66d;4IT4c0LXG==>H9UbKNTb6.)
N1XSV&TNSIg\9,UdVbe.YXaf#cUSdb:6KB<[JB8C5T483407@4D2<(dDN31Nad9[
?b)8/OVgT3NF36/S9FHEZF5#41O;@56aWF(KQEgCRCMO.RbOK000\>fCb>&(KO>0
=K;QI+\20Qbb+[>#8JVbfN1HG_E>7dF5Oa>dLIc>ZMNgY/fd5]cMf8@@g@VA/8JJ
J9MRO\G3\/_20-5ZE.=NcIWGKI&B94MN2AJ\2[Q01UH^F:N-D#GIMgdE\[IQ[?3P
HAGW1Z[FV+7^g&N;])RS,X1HZN],18@1C0X:F\a(4P(>@A,E)?-T/7fUWBKcEFJM
HS8<6Z)L),1OH_B6:V4VZQ<\b8N+Zf>\c&+#,K?N3_.ZNF#A1dS<9A7?(4[_^+CP
N+eH1]1E)e@#MDTJ:O<>cJ7H<+79.2\XL8bUSTJ>4bQ?9W)@=8AG1L/S&b.148><
0c__e21@4BMC&7X2;,:_K[=4ZU&I/4]-U7=[1G?:G5bV)Z-V8<=V_.)[-a-6G@Q_
G&V0C1]6Y<g^8/f^)Y1RGIEZ,d:1B_5[SA>ObM#d:4K?0N&=+-O;&C?D(bH]IXa:
MU:OYB(:(2ZfRBYH9?L,5,I&ERBMG0(&0KTa4D<]A9^H&:=94e5bX.dQgc[H<?V4
g?bKaJERR5KDge0T8OLA(-1.UPX7bTQNbH[>>>@d=(.91(#@K5+IG-FBWE+],)Ue
JQaKU-3-d2:GTX+\g11J)F,#))7))aLH)fA4aQ/Z6fXVf9>U:77EC/596]aL>)?;
]^W7aU8e@S#2^NT#;-_cM,-8N5b#P6VGJ<EZI3f[/[W3M@E^88)UYgf?IY/X;OZ#
eV+M]1Z@[9@LfPDA)bOM;(K2XeeW5Tf]=GU:d#?;e9,6g85.G=PAW@T6SR9JFgQK
a8<7A,=&3g6W^.K,AUKOEIF6><[09_YX+F/IX.8\IT8[6DX?7@0\&S^Q=0gf6ZJN
eM3RI:ZS.#\.+7(cFD):&2QXc[B4aV6&#9-&NU#[6Te8TO=>DC&R7Reb/0@6OF[-
N930DJ@TbWQPLI_f_=X\V?7JJMPeU3616Rd\J\0P-=,708Yg6=L6C/>BcR=+bE(P
,gCaFK-R2IOA(XI8>I3.LBQ+@O>-KQJ3-(V(BJ]/U.;+@FaM;^4P0W+J\FW<@Q6I
\EU)((J7a56\@a8cCGMdP[D^1,4X#E0R417[&\.e_FR=c3.d2T)fGT]EdPG>B_,+
F_O,K2=-IO1]aAC169Q)#H-=B<b9Dd7RXL[gF?QIe>]^DK@-+b9-/ANGMZ9CaM\S
5ZG&&KIIQJ8<5I6Ze7dVd\/[a_.7Y7O-/aFdd4Ve#9dANRD@J1Z#\-H\)QGDc2>J
dAf^+8/BR11+0_bNZ:.K]Ha=JWG(R+B7M@R2[[9_;.,X/\O#.@<H_5/#W6H<#9Ha
3_@)0G+-];]8UX@6<d\2@LQaRQ]@PZ97=&>?Aa<8dQ/d]-#[6XC@:)_BWWL6e?_Q
<HZ=8e_P/cS=G2EXQB#g4,TWS1>d6\ad#50S7>bfX;4R5_-7&=0a1GfV(_UWLJ8W
A^W7P@I>?/b:+4\<Ba82W6TZ:fG1\JH-5.YA5JJg,9M<\D01N1;-VZ0bLVC].X#7
+c]-J)YQ--(M0_ORPZ3(=4g0IBWNWT.@#.eWA[@N#IXP#e^3:/SZ;L2:)])a\36\
Y3@BLJ,AcJNW1IK^cYRA3K[;I1/\-6ZK38&1ZNW-,J;U<F^-OfVXBN67gK?(<\FK
1=WPe]+N4f3b\SRQ\FJZE/Y]5/W);R;X+T[TE2I?a)R#&5_C+1&M1PWYICEMW2(.
WP>K^KLIK6?aWL6>J&R+e)CRYU^IAXZI]CCC<gPgEF:]7M.(fV/Ud(&?/&0fR-S=
D4.&L<g=U\EK#(2M-/(34dG4THF^K#-35)Eg<V(PbcOZ6T/;G-D8VbPWg0>YVZ90
IZbA9,bJM,-986KS@R9O:YS5/>ZZ&<-\SMHdBMR>,W-L7.cfMZT0)T@P7Wd2c965
5Q3^AP2Q&H4N.V&;MIX3SVf#gXH5.:6Z^SNB9;]NEAFV6WZ&HJCT=>_Dg;KMY4:6
<&U2Z?WVKVXZUIeL0^GME_@:0HgF(Ub^TM<E>:K9U4OIN?=?O=UP?bXQFX_5(QB(
UbGX,R>Z9YA/FFB,g)1A.LFY7MV[Lf;X,7PS3W\f>#LRIV\cJ4f-B^gaB;OQ28DT
GXDQ,85;0D>V7=YM<\X[_E/^JbK<N9<a/78PXeAM:(KI)2dV5eZJJ-,8TT,bN.6P
3+@ZW<VGB@E6#O#9g;>gE.aME11fe.ABH3GJ&c:4Wg35M09FN0F,1_DE_</a5I]T
OgQ9>R3Ig_)g9E^2EgcH^INb(VX1>a+85VEe9Z=2T/C)R);f=L;L=7T#bM4LVDD3
FOA2+0E\_I9EIg@WGC2:U9XB((,/Jc2E6N6(3\A@+2(000ca>E>;f=g;-)-MGCMK
^,Y6_2ER:2cCNJ/fO3b5YORB,:JXFEGR.IP20a?2+H3YbXK4YN+HfDZK6VVCB[a@
-8_Y7WG[J#:XZ@#dQ)\B(=:@e3>(40@>PgV=/V1(9V#gA>PHcCDd[+VG.=VaE?IY
@GJ4R^(6PDT+)[]+==fS]W))#,e\Y_=A;OYQI0g-^>&T:E_.7SFd@:Q,@3=&Y:@X
gUH5V:Y;,0=G#5FE-KZGX?M?1g)_8UN@=fJ);&;M0L(\\CDc7(0I05AbX^YT\;2W
)PbE:0[b&S6.7&NRe/Yd90\M2PU?:-2?V5Z8aSga^F<@4.(O^EPE)YTH;DZY3Z,a
0]I5<K]&VdA=C/C2MZ]Zc0@T]N,W6^3b[,Y+d)1T7(U(e0(A1Xb61-VbQ?MQT5f]
fN<.S_3G=L8+^HVJ^WHT<683R=\K[FA>c&0U(DHH@,9,#<ZLcgG2f91#1B?N2T-E
aCX)Q2H]KT=gSWY4Bc=([I4X(<GQHC1PcZPK,4?J&T=>Jd=,(O7B]f#PKV-YaEgQ
,G]H1Y<Ob:82g(WeNA2Nc008_@_UZd@,GLE^cfaJ8M@_MZ7VM#]-ADD17R+JT5KS
+4#AaOTI^d0&D7KQ9f_K,2:(11&F\eS5&@YJ;R5CUV=L2BA)K\DV72XcPPL7_g-c
Xaeg2MaRM/4?H@=PHgf>e?Q[==a6(=4D:^C+cIV?QTYR4?-->>]&)f08fSO4EET=
(S/>+^)cF=)\Z7d(]U=#)A_Z7fNS95EaCRRT&)7e@)\TT;/+<-Q)/gS2,Xd@YfH3
Ua;.GIP7b[bg3#Z_D\:NOb8HX7c)J@4NJM@H)5S]eN;:Y]-TCWY-RO\7+0VJ65<W
///DZ([FX;X810>^+AeMN3=S^JQ8/33=gcVWab^=F^2Fg(60PX;@\Q=W0Yc]L[Hf
,f(U@ZJAX-MQ<?PL&SAGd3EdTS?)^1dO@=]75SbVO-D1/A,1fdC>31e\@EI1@HX2
#bga3?[6_.;Fg@^_+(.cT[.-^V.6gZV8OR>aNe@08cP<D-O\VX,1I?OS4MaL7]C-
^e:)V8+X5VeOgY2BTT5C8Q4X^C\L[_<\6;5C@3cX3US<g9:Q9YGK(E(J&W.8+cTO
;g]Od78;47<L8P;EDe]Je(NV8Fc#Y;4.0Wb8;H5/8MU;N?(._JUK0cEaDR//Q#.4
:1LJYOVg74A+b)g(WDW)KaML^Ob\.Z80f^XHUV6A9?(^6e;UI2<3DPM38JH6dba1
]bT\aZ(RF;#3Z,fYVG##,?d]ZJeA\DN8B&,fT\MIS4F_--9GY4UD#?C>7#f/7&NI
?4QG&\_=V>eW<c2:/G@RZ3#Pd(;c?8Sb\)A3,1.:,>MM3.6MbAZc4_XCQJ74V2ND
2A)/,6_=&OaIeJ^(WH(^6d8HE[)[WLPG]:DPCVC2B\geEN6+,VB:JA>L\]\/JV.E
0:429D/8WKX;aM-e+W<F18(ME<H&VBK-8.B1</).7EU5Cf:d+01Y63Z/c?b8Ie)+
\+_cS?ZF&U=JX3e\LY)P-H(?(/#T3B1<K;4:>9[=0#C13db&AdC8Ng;NK_V?,&27
g.AQGb7A?E(>D4YdDD>=cN#d[:7\X7MJMVRD4@PZVgI-Vc.QYSA1aLcc+B5,0?aT
eVaA/;#G/Qd87aE><e2T.WaK+D2L+])X;6V3)\W2>[Sa9a-Rg_G;TPHg^?aN=:>_
TU1\YM[#aX=<2\7g360c0IAd-?<O@0e6^[1,@,7S3Ge?NI@8JF;K+@efa1e)TV3I
=WKW8aS&b?g=20IPKH]@IfUR\2c1K4S#2&PA(:-9&+Qeb=0H70UXU;0c[bF>5E51
U5JHg=:+)3WG8GdO?KV]WAT43=TA;\8YG&HPNbZ6a#PO49D0+@IB&TAO1X[_41I0
fJ=bI,Qa/98Bee;LSW&(4WQG.O5Nb0QTQ462PX<+HXIT5(6@e4c]J#^(<9(a(X0=
L_FKN5(c+V@@W)OLXQ]gFTWVDb;T8Q(R\Z3=2K.fQ-Q=Dd+f^/VbQ2A54Q;-:d=;
0F0SORO]6PMX+E#GE@H<aO(;\N@C]O)3\;@.E:[N(6A],A0@_bCI5T-@eNKL0SUT
J0-1YPBA@G7>IA>Xf1PR&#OI<dLOfaZ9#F((7g&EOLb)H1V0dS=C=_K@<8KC@^70
JQSEKRI1]R7Gf^1_.RW:JN-\Gb]-Of#PWRT0S8a1-E7JUcYe6HR=LKdRVFa+:^;V
CV/aage:1L-+[R?NO,b1Nd>>6G::5FO[=)7]MfbBB2KOb;&2g#5YK6VY?KIH88S(
8VE]3gQW(X\HZ8OB3\II[9TDgO?4DI]K:9J=E)//(3e2DD?)&&C(9PYYW&OGeNON
#JBX)V#8\K]L#>@3=A<0-J4X&]:d9O8WLZO^A8MUb7N_[TCF-GU><(<:DE2V2eL8
:E^V[LL,\(E9HSSdK/YgWFVDMW)-7fg99Wa1DC/EXc25PN84=33#F#-B:S-Yd<++
8T4eOIUJN.]S2H3T(D:DX1H<HX[3BWF1D4GO;KaM4YWXF@<SQcd5(d<YGYSK3TQb
]SQ:B+),#a.:U4=GN]XX@E1+P:/TY:gK?(207fX6=34]55E0@S.I=HNDV.KNGVA5
J66-^OW]gBECU@?+O:36TJI_ObDd=/2#M:dZ:G3PJ_I\]CaG;O#X?FBWD&Te2,OY
JDIB6F8E#XX7f(=)1c4+K/b,36R^e@[7/^2YD[&FWFdQ+</E+75gE=QMRbOTg/&@
ZVVafY?4&G#,EdN0W[B2VU0JW)e&@2eV1D-(6H7&AB@S.KC(L9);5/,<(3F1&XPI
/e)&D2=D@Q@agOgB8HG>(_+G.[+5g;beG.Z1cCQSQcRJ=\29:g2SggH&B4XJ15D_
16PNcD&^_<E=&(=14=O^_XC4Ge6\0?DQf^#(^@bE;4F,-[d6^NBHcGe((NZWe+M0
#<.),Q=E\)9&#:OW(=K;CC90IELX>gYZWUa8bC<ED9)?PEaF4d82/67J(R.I]<#1
#I/H>U-\@d5J5U2]RL#9bcK<T,<]B@=WB,C(<C</(Y@-M7UOQFCg8>bCKB\LTQYL
RAZ7FZ;/7>/d<+d@+eV=#[S#7^D0YU]dR6NRE36(]\P_;5MHYV)F6@=,L#BI>_ZB
)Rc:(=WVe/Y0;[<\bZg6D5>G;)<19+NT&];f2VAI<=LV+T=gcHK4)[EOaOXeWfU-
<AL1S8eOGeG\&XX>d@:a(&_M[bd=XZU&-_Y:YB9:Md=TTL>CVDXV<P,UW2?,VP<\
ER=;;f/-FR)7_&-e63J7GdEM,f;S/MGY0+Y7XVg<Og=/7#aGX-YMO##T;NaH_g+>
9DUZ0Lde7(3[J7E0[f=2:Ie/7dYM=[QBc-+>_Bg+NG]):8]5WgBUY#=RbJG^H5Na
O(&GSEENA@^e.I+P50-8+3_H/>^2Tc)OXHab,,]7GZZX)dd7X2cfH,?<]d\]=W0)
P3TF=5DI:?Og_=<6QDU8A]g^<M#c5_RT[OdgK9W/L)H.S/(DTSI9:T?Jd<=(S[d<
C0<[O(4TOBX3)^76E1_d4_MJQ:?(?]Wf>D;9V]JEYC?,PMb;X3AIB/R<dI6d3Ed[
E;J#LP5T<FP?-WPZCSbA2GCK@d(BF5&FcEZF-SIZaEJ?FG(OYX1Ka,AZ0a;.T<7)
+bbVd5^.U?FOT-Z#15L5Jb74;&+>F1NKYNFA_,aOaR#a]3_NY&J,0Z[P1],SW/(V
T2?>S6]\):\3EOTK3-1ZALR_QI7TTBBA1-/7H1DeV<Q204/#E7D?X;6-235+X&R9
UJP)a&6Tb0YcSFK6VX63ee_A[1P=d)TBH<A6B>XCf=K(TPE>S<Qd+@&Z0NCe1;@K
10eH/7,^VIUA@<6_C3g_PG7c3#;@]4GFa0b&Kc@eAWMQ\K4-bOEFb^6;]eQNZ1Og
.Y+dXXM;S\g^#fAJ:]TP2(1G^#@[(6Wg^#;G6;AV:M=]&^X;^g7+GYHJC=K^FQU=
<U1@^6X/A9^;\VZQ36A@99+G6:?PM)_VJfa8ad+:0<UBUb4;MNg#Z@Mg-&ANT-IS
-^>f=YeA@W#UIaDa/PUfB_>L8>[P_T\gZI2cb73a@U:K^_BJT@Ag7#IFU2@_3dD4
RKg>8[6KaD(f>4KL4?[I,_9f(Z+7BTHH9MQ_XMWZP/0a<cV<^:JT/,O1e?+LU8OA
T#I,,T#1W=7f.CYa_2F;1I:gI\)3,Ig6MS=,3AFMA6M\f&@-AX:@.TEH=CZ[ND7A
Y#BQ44.FC>8D<PZZC.dS8e\<WgA=.+UIf(cbO:,,VbCJ/,C=M8SNc;/ZTK+D+UOB
b311@)LD]Mdd;U&=]YE9WFe::?6]_(.2=]e_(:QgYVV2X4F]:K;0M-#3@NLaSC4F
P9>LgPF]&59c-<db)#X5S+X@59X4a^SP7=e6-1BYHA;(;HG,B^7>#c5P0-P=;8dT
^B6EL9;A,KSCADM?D5,JV/SMO,KRW)D,X-bA_IbNU\dC5bSV+G9G_=8X-/.>._^2
g^g.[9dJUEEe+S]We=#3JCOFXN.0T>.#(0-9,b0cG7,^L7H:gMIV^a]UI0/8M^2B
N_.5\_^NV?K9[)F/Fd@H\B9Pc:RM+gX=D0Q75\+3Oc<==DBF1b9DXcQ8LTU8.,?<
9O7L/6S^ROB?94GK#S_J#0GcLKSWeK1b6TT7_7;]4d=71_V>f#9-^b#:0(g3b2,U
MN)0]K\[TXJCN)+,[Y/>=03EAcR4E#M70<X]U>(HOL6YOSLE#<6X,Ka-UA]WC[3M
WLc=B6]\1g=7c+@5V#W/2P?,9=DIC8VgWg@>2/1;_>B8f#^,-E?DP4_JedFZ/\TI
-GPSaBB^Y&M++cUcJ0PNR+;[0+-+,8aA#D8M6K5dbc6>.a)C38Z,=d6Y6WfD1<>V
.@RKY4SD[,87=g;]QHTHeB;4]?_cD4O):JW47X2d1IG[X>2]La/=?M@dRHbQX2AY
-;:eYQJ&K=B?f?5>^:(?BN2V?[?a[2A2:BLbU<XVW[bB1cZ/MD_3N(3c#?(X0:ML
f]OP/S2G;[;V<FL^58(C.:XEDO_GQ7)61EFU<1\C@KeV&2gf=7Jfb5?7FS.Rf:1.
ZYd9#W3U8S3[->=8AdD?7[?CEW6eaF:S-0VAF6U0P[#IK=Y64[@W]9KQa2F6CBGd
>gSCXZ]_4OYOg=N4OZ93e(&+VH/)5Q;R7gSJNN3JC2:SCe6^0VN5EYV;[F1;X-^@
87fGdA1ce=fHQE7Y/_L>^5+eO#M>e^6@OcG-8].Me&7K+B@/K6C#g,dD#3L,TgF_
QXPPfd>RYC0dLD6&3F]K.ZI2YJ23F:UK>;c,7ZeY/_:=6ec:]Hg?c9&;?MVK@+Z8
>#6KF-0Z.@AK.PLRd26TaV_GDDaFa)FLL\Q\#b)?4L46M.Q@=/-Y_La[_+JSN@2&
>-9]:38<W+#QLR5(=#bRb+4NJcg;WN<cL/XHb#IP(O=_bNd??BbS.W<6bO-MO)c)
<1)1C3eD^LfIF?VW3>g+f49^Z4<MKT/KQ>\9+MXF\#Z<f#T]WdISXga\O\c]V?J>
(5bZX0IZQddd7bUZB\=_X[K/K8IX&Z52)#f@F]G56+C.g?dBE_,H:Z/+RO(>E^.L
2/=)&TdBSC:NBPb<2F+;1bf>XXC#D\dJ\H;YW+,PZ_SeQYLG;R#(\S#_<QV\GKKa
)8P;RVN0WGdF2baY;SOb778B4;,=?U1CMM5\Y,?a0a.C5O:8K;6VOI\38D(C_bNg
1?6Ge:&T[N:LVJW@ecK-#(g5.aI+<I1,)F@P5Rd.?\FD7&RD<8675^NbZW[@#ef@
@-PRD&cUGYfN\cd:=J285AMR4#cB(U454WJAf;ba^)RQZ\2d#EVXd3Jf8KN_[:PN
K2=c&57E(XI(3DLa8LD-T_SBO-STJO>18.Q,MS&GJATE2)G>Ha,C2LW]d5IYU@N)
IB5a0QB\:@=[][NR56I2&@+0ZE:S8PPXgK7aN4OaG[c6@4Nd@P8KF,8^N-LZL-Z-
B\=<+QC@fR+U>FH@V4H&;IIF66RJLcVG<?aaDY6W+-+LV3[9bTg3e2XWY#XG7H=E
^-#a@8T_Y0_\2aGHYHI&D+.7(PI495J(\]=9N3Jg7gF9/5SNDce5Sb\gE&?/ad6+
@]XB\:+<ZONJ:O;e1(Z\6W,CURL.S7g<G\Tgf1/5L]RG4#[F2LTM6TP9:e@8^5^T
:(5&^2gF<IgI[74=11/76S)YR7(A^=HX(D]:ERJ)<E;+beK5^3#(fH(-.#@0)/c=
^GfAWA4V>BR4CQJ@]QRcKZR(HGF8:[05ZJ4>2?DPAR+UHP;D<&gTD_9&RL.(EE64
eO)/cfFdEe(Z)+CZK(Q1AZI6,LR+5]Z\=MD=4dXe0=A0^^M:H9=IG?Nd+_d&E.L(
[CE)-3S36T_W5#?98GY.\d+g[MBJ.B9^A0:+066-VfL\NZ:A/SdcD9W:4^5EW#1/
(^:<[\b\=I:a4b(fbNb;]-3P6KbUM72P?=0g2DJM\2(#HG(:0]I?dT>J#07ME6fd
:+GXGV]e3Yd#e9/gFJ#P#FTER=)S9\54D9XI(6V#\77/d@+e^#XA9TGR5f8..J+1
,RcPA(<M1]^4[C.BU?,93OY@VgN+_WP\_e,/I6FQV2U@WOPB7;Gg2e?FgC\:g-T7
/Y@0fBaeOLa4<-;C]9VJ3E^B6(HAGCJd,eALSZPaH,=0a4WEdE)>)#WM;A<g@94f
ECW<8]#;;-7+ZBUI_PO:QbK(A?WQ#_;-2OHT2P7Qg_3EZO]85X[;M,DD+86^M>A0
.6B]VCXG@Pf[0VZeI5fZ-IAa,:8Xd#\g(eC4G=TYd_d/P8:;E+J)Ve@&4#DWDP[R
e;H2;[04],PYJ=E8;+&5CI^>BMHM@XeceP)#XaZ<HH:\(P&V3[N760.6M;SRNac?
V)CR.6\DL9&7L:-,ERBU=SG,E>.:>749,CAD_-0]FOZLRe-9.=QGXE/2D/eC)3e+
5=d]E1cBT#83Fd9WDEW/e2N1=QQ[GCc]R,0fe[RQH\-5.1+0&81,TISX=7E,^_\P
0+XHfg7b@g1U1FbCH<0QLPg\5.463>/F1M^XK._O?JYP3V7Y4=.JW5^FK>57=9&Y
=1;VI7^(aaFRBEWIV8.LB:22D;eE<]>a;I:N<@2E)MS?EZdDaMA9,-g3IePJ&1:G
2gcOU2FcY>#eE=G)74_=2]F(L;D720+cERPaadVL)1gYQ,f4Q2.I?>:Z4BYcUK?[
+P<L:MWZ[QGOIG)T7N65)dfM\e--/(6,9+?>V>^12HYO@^OPN&90+\U0W;T#-_IK
/_=T?8@FM^Nc\-VFcU4DEBf:DXf)RQCcZO(K0E:IZ0b#dVB#:=cZCe]>TX^dM5BR
2PXY83;Jc<3QH&5;=Y.a.&eg_NZ5Y1U8GDeZA/C+N<0XDaWdE=A2ScXCBS8=JAF9
,M#KROc=f/X;F6:VE/Z.N]gG8dAR0\H&N5_UaF=M&+;;EV_]7MOg];6R2(7d9>LH
SSM&?B:,PCNU4P;OY[GG_25Q@9U5#2FX^@NB0:B1XCcU4Z(bL:f>1dNabJ\8b39X
Sad6f]>W844WM_0-UO)c/_L)DAgP0aaT_C68099ZWCNMN;COY/7(R)ZP&CJ37\I9
V+e)6SA)]6UH+2N9N-]7:1;#OL_50^[+5&KD?V,#NQP8A98RIUQ;Rf=9\YW>f9PY
aIJQNE,3T_<9HM=BQG:(Z:]KD_FbLeM61:dM]8NLF/IT^K:8Z]A8ZI^J9)PTc#C-
77=[#g&8RN+g0&cPTaNP5=dEfFOQS5M51<.+_#VU>QI60J#c<;QNGL@BHZ8:,>(0
Q.7M;;WF7VK2\FDF8EP;b0//J<48RRg8>c8[aMJZJ.12:2Ia3M#55-D0d_6M#;.8
WO,:UZ]9+VSJc1g[XKTW6LbNFI^DX/TY@KA.3gaKPGVSJ=d/]#ZSUV)-+Q.Q#U:Q
S_FVAcR7>;95g]D@ca9<BC7f>^+0UDN6NYg?5224,PZXC[3\),:=0.9fRN^TZT[[
PX4P90&()?Q\?Ia@bJR/5Xa[D31VIS,I<<[D[gITRT#\6e)1-&U_#0D)H/6OV\Qe
A5U/)d-4YMBeHKH+MC_DfIOZ:MPN#8SYG\NU-R8<;H9eDPdV38Qb9B0OKBgC?&P,
^K=VF.P_[e4/B3,E;0JgZ[A?L:.#MGRa>RN#B#f//B2gZL6L;D>_MT,8Tf?X]59/
gKPJ[;3Y9;+\79g+D1#Y4#HN<g2\Xd\>e(YGR><MZW:^&0R,P<+FB30M(J\64TMc
+5685YYICOX052c=9g<9(M6beMWFg0fN-e+_=R[.33V35R[7URfX;,9EXT3?D\0O
GTS1HJO0Mb\BdTJIa0E4WSTg;HFJ=7-^?HW3S+NQ]DUL6)_F[eF.[cIJ1/=)=7)-
TWa\CTV)?b)+gW&?T.UIcaNT@_P08+IO#(PFg>8O[=KHKZ-29,H,gdT4R#;8G[RF
IVP&6:f:.aX9^UYK4X=MH=03JR098TWR]fN&8Y:MP:?d5TTSY/#KA=A7#RQI(2+c
8de>UESgQJ+J0):-5+?0aK;T,&PWGOUeI0&CKa]GFE?2\-a]<:Wf:fZd=5g.cKN0
AOUHN+_HN/)6@IT_8]d&5E\.[/;MJ:O36D4^T)[F9I8D4&@?Qf+(c\G)9-3a)GA+
OCf[A@>5O4::.[Ec6FC2dS8dO9eQ)S-0-\NPI63+054-(3G.92?G<0OR<5Dc:2MY
7@FDad/Kb#,9MF@RG[]La_d#RY?O)]60X3X#7D]_.3KNA&SO>;1^,4_=KZ8#EDUU
?Z(82G:?0P.WB3dE5b>L>;S0SCYX]5N2&Xa@V410;ZdV>L+M?d44_&((4.VMBO[Q
XbQX/d@-G.)>aYR9I:=B\96SQD9E]A=F(W#@T365e1;8BEI1V#bP-D+2+Z4[C7VF
I^15/EC3L:;dfGO2b((B:TQFeEB-IO&HY:U.cEd;[3II^E0(<N[c&FI800XY.VE[
,JgJ^FOY]#.I]?dBAGfB1UC<G+<8d)0b:c6),+-PLeB1@A8d);-dW-DbD7=Pc;VK
EZ;BKCc]><+I[5QU?Z?O]._6#BPC_@P^6e\TL[G_c2Dc\4Q.^3L/FSV_KFC(fF7(
ZAeJ;XN_WI/eMHPD4&OO)+C4Z7#?3Yg3aU_1Ff7DD9c(L[E8-C&X&XF)/3:[dALI
G1_cL_A_[:L5Jd/Q5Z4b\H##L\\WB+10=HRV6LRSX/H(EN>]@CL:b^e0OM<J<+EZ
04-I1JReE8L7)RW2Tf-8bBSA;1\b,G_]9Y7O6Kb<g.++C=@#O0;cgcJ)+cYW5Cbf
2N\\9IU?F<90Td#Se#]]2(I;@M@^FcEJ--N)IY@E#AIdTN1>F=TYgFTDF[<8.EfA
/0?>d<Z0,3H/S_9D=>LK3>7<NG48EU60[W9;;J4R^9/-a,K1^ENb0SAR\.F-ZB8c
AKG>/c/+=,J>487fZb5^SR#<7>:7&2ZM[EGe[3+P_3TJcU041bDHV0DJU>ET&)Ag
?>Cd6fXW6ZF,SOH)F3&K+TKc,N.S&de,LUSV2T=PJ\0L00+>^JFV;]@S[^-&:ETF
7]eEHX\bWM+0;Z2,,-fHM#]/L>V]YQP>3JMY@f-BF:8K,C_A#QL_)0(#R>13Ne2_
eU?VHHMF1eDW950AA(^bAZfI[+R.+J(K@edV&HSS9QKGa)QRY9/Z_X@>]<bZ,H6D
2LFP-:1b,6+N:&1D/[T/C>29L4Q4QC3[412N>=RP)-<YDL_>;@-N2FNQeG9F+:=P
.cY\]=8[YG),C[]VgM;c;?C5@+1U777_,\dfNJHWK2-^S>:0Q8LJc;A2)-2)ZR(_
.J?e@2c#5]RHQW5YA)WS^A>A#=#LGED&?Gb->DdGde\V+?X#5/.A[:3ab>8N<S/_
cfY=dU.OY?-La+WI28>\?+Z:@)U8)8SGV)b,@Q+:S6c@WE0N49X@0(X?a7cD]=8C
faD3>J@_VEYEPT-(Xd(e>[E<T=HD=>#E0_7)(G2e2W)a;YZ(4:eXPPT@XA74Qc5G
N]eP0<E14H>B:=[@;RNL-eN#>37-J5JDD>&6UG<<aE<1VQICUXJ<e)/C_.K=#G(I
H)&CC+2NO?_f6Q]g0^L)TVGM[-BN7WLE]-ZOW2)HORgD#f);eG/)GQf^[D.+IKYH
^.?XO.CQY96L]b[M#K(0ba]8d])]1/]fB99G<HTecdKIL/]:,3?82ceXHQg0\6PA
BZEQ/4@ITBI6cRTF=9Q@;e,N+W44A0J>gBYd.:eeTO&;JCS[C#9_2E97P3OPRgVS
BON@ZDJa836J,I(aLfUO0-JI:Na@(]G,Q.&7<gd8H\JV0BXAUP7QHC8/U<A;PcRQ
?.E720^NVK/#S\?U^5U8JTfYCdaYa0Y6e_8HF1WS@2@+&#--P_fe_F2ULS0AP_8.
6+:V/O_FSKa/+<613P7)4H0X1;Y23AYUb4a&GC#(RMBU(JbCXK6MD<cSP023efJN
>^YTL?/=f&TY?d6LACH?F&>0b5-=0UHYDQb00[NN5ScVJ[G<S;]4R[b]94T_A\5<
TY2<6=&?dT_XW<R,RH5e/:YMC62Zg3KJ\R?^G7AAES4]ab&QbK^5WCNG_CNJBgaB
)f,f/#,-GGY,NLJ9[FM9,TZd9BI+Fc^4OH]OQe6AOfFV(Q?5(@NKcDccXG;Ja#;?
>aHDU?c;YK^7g.PMVY[1/\JQ;U]c++[2:<7,fN6U?_\].:@-SQI;EW1FLbQ04XS.
UKCb4e.9>?aE5^c#[LCa@M@=^A99c],9(0,7SIPD7LYSQ]>-K=/=0[c=/H=U38<g
^VYNV15aFI)L:=1b7FABX92OMLJQ589N:91:YTE?7?^1TELcafVBBBA^UC3BX0<;
<DNf>4=;begOf-RJSMKT1M4FO)^;]WY_?F7XPVJ,[>QAdKe[f7MKQ:=-:V^VB_G?
Ae0N)EF?;7X[82,9CaPI(3aaPGH/aG\O,MPe/6d412HM=>-5/45A)ZNdQP@ee-;7
+.6,U/gK84K]G?[)RXXH06293L,[NRPWa?JeLF74VMQ9-14FQR)26ec5A[_1QRC^
44+#L:CB-eL49>?];42<B]#T9=NW?ebZ=d#LL,9P@Q_YKIWYD?cP(3U.670D?fHT
?B3PLX4P&H__U8#[e09a]M(C^5J1S9:FAc;>a8A#7/K8<ODV/:)O;(RY/]8TZZ;d
GeHC7?\59\\YGZ&^HK]K1cG>JLO,\^@OO)Lc9V>F7RWTP]baY@;,AD3V#PD&f2-K
L=0(QOZ-R,/]^B3_L[-BJOdJKD4g4RP5Q3H[S.DARZ<-=D+_=@Q18&^L;RDd:IHg
>79A_<[VbW;B.Z=e.=O4b/7c4)e5e(e9)BI5c#?4GCUY&HV-]2Z@9^3?:Z]IgL#I
a4X29_VC7H]KHg,O9(2f-Gd6><.[9=SHUBH@UQIE8=H@XEW/J?BZP<7\WL:M&JM2
dEZHVcKUQ<g=[&-985L(43E,,,;8V6J<\KN2TUd7@GfGGE3O/)>2S/78g=A;J5S]
:K#=J2E+;Z1ZE&J&g<(Jaa9\VJ5\>4,JM:.)?:<\K8K3^^(V:6g>SgM9QaZ+(I&M
EGUCT6]Y&:AFbYHBU::+B?ASXd+I)I]2^SDC>_O\Y?QFY2T/A0^2.=I^O-0+c;UZ
T2,GVeS+I]4&NT]Q(>V4[57Z3X7K^B@/CU#VPCKVd&8:&3ASAB73b9#@@f\C0G._
NUF)P@8NdK1U1K<+0D3e-5eKJ\AaY]TV+1(2HG^Bg]b1,[Fd>?2#c7TO<96A_-/,
W,bRZGXY1VPaa5Y<5SFEE[00Nf(ODg--J=gb(aFIH)Ib#2MU@b7.OSWZSYOXRC8F
:a17_R5W]Y>Z>((X+V+XJIJ8JGfWF;YO/&=YWE-1LC]b9ZV56SgR?e+L8,L7VAF;
2]97:#U>fb5P,gH1AcTV/)bcX)Ig0U@M/PPX6NVX2327:^L#H,O:Z6[,BPV1;6=C
Z=U2DP[W2\MA,VRW<==dW^_TBOf3X&YK0OS/_<DgIN3(@]dIFc6He7GQ;6RVe_8b
d.\W.6ZSAEA.C#0U9L,T?O,G)fS57\>>H^^6P]Z52946T[,Q[+S,UOX7EL]W+_f;
(>AcJb8IR)CI?]UG3C.(]JFUf3gK/&Z.:a0SW9c^1_G6Z@OM7E/V]_N(SBSd9S?B
cd)f(1>2G8CW>S#O#8]9K<L]W0UI_.JUQBQWN1@GT^,3PNER9dEDBGc.1aXbPCPZ
:)eMX./\R@D2&IJ#-6f;_0\L-0\KARacdQ>Cg#OBBXf+KEbDdJd6GA+]A^C#Z@@.
C?GV.O5-KYH2#9g,TF\#=6fB/DT16N<,FQ=:NED_6LLRZRQKYB5c@-X^;<K;adYT
c7fHbIF&#^@<MR.-X.e:W(&7Y]1,HC\/1/K2-JEO]08R>]]@gW0>,M51Kc[]^.#@
/cgfTWe5J-CT_HGX#P-PT,;2:VXfDFPJ3\HLLd6OAYfS6&]a;T=1I@A(NTY6aE37
ZWHD(&\;fL-@PWe+X&=/],4a+UP^7dQJP2K\-7?NC,3DK;BP;W/WegUcF+APHGQW
C6.>4TPOK:=HfH#K[4P@9V(J3<.7W^(=a4N8A>V/JRZ9a(0O#QYeHLNHRSJ(OE)d
=XfQE9DP7L([5_[e(<?,L-GQ4>QD1=a]>95:OEPNQgY4EYMVICV,bEK>V.ES=b^a
.]W@LK@dd&TQ(>W(QQ0d07AYJ8IM],>CR^gRBMUS5dE1YcJ/;Q2C3RYIEG;UO@:V
&9XWHRg4&a0f04YM6.+W24X?XBN?BK1b+Ye.W@Ce<E2XL=4ASFY5COJ_>g2\/J>R
M9YH#bF7NJGJ;.7BcVQ9d]Td?c8gcL#U95I;5/^(MKU-BS,\7>cA>7+\17[PW+EK
gRF1@USIFV\;YIUVPS(^A/&>fW,Te>_>:.=>57N7Y=T#Q]eb\2^=--PWKRDKMYLO
)RW>YI,3G95[TY[2)a5?P()RcAZ]2.1E^>e--W[#/EL<]b?UAO=e?V)36a<M.KN9
024M#?eYW03K;[AJ_BI7/954Z#:-=12EX4cWe_I@g,fB2C2RSJ;\\g#>T>(@5&U:
T]aGA(WC(,I[cXH;GL+QS4WHA+,\+@fT>0?3gM>0gNO5U-PA0PZI@;RcH?]=d(@9
FZbG4ebAf0@d?&W-ZT6,2D[ESb3^^27G_:dUUEaJC;_T42cG@VYCfXcSZ?Zb&E]S
]:X4g;&9T/I^USK/8@:XEXF\Ib.EQ3Za<KP;@BX=/\F[.#@1CI&&F#J^6gA89aKT
CdOYMKD6Ge_A[(7#7PYMP3PJ2AXK71(U;/HMF>671\,E@[[\UdFXc9f==3W7K9=J
)E05d)E6JQS<AELZ])6K]>N,YW+4EHH#@C)\=_I>d>F;TCYI[K>ON16.gYW+L9.H
N7Ia/C(_)ZAP[f=Z35\88B@?E,LD0EA=L[;E)gPTgY]IX/Wa&NX^]OW\8A\^NOTT
FT2_47fBC+acAcIRXg;7:d9;f</dJN?81BbYZI:1eS@MLc]4L0T,0E.GO5(SDQ6M
8Q>EQ,<X7.P5J/aLKT6<dYJHK>cR@UA.:#1-)NWR-M/R0&2#[-N<(^d&12f^3Y3#
P&KEHJNCJ_W2J_L9X2ZK1^GCRL4P<RBbAM#.OU:f:QKHYg=DFLFR^D6b@f^IR_BW
2M?&<CJ###;O:G9cg1+L6(^b_)DaW3ZQ;,L\#[+J65cWLICU#B=>##IQeXW\K2BN
[6&]NLCO3_O7E,L<)45+,>N_7[cYTH;PVdeX5W>I<,/6+#:[(f3?.0^A0f\#AX57
=dG4W-:MBIZRF<T-FW.DGL5IQBY:2Q[#.9;8IO5#+&8_;+27@7Y1b[\(DdWcCH.J
?a]#T^a:[:S5V?>C-aBX0YTJ1>31=(98baV/=OH;8[#?>We,7?8c&#cRV<8OM2Hc
[KBQZ;d;\T6<)H/MR&]GCIdE4::Y8HGE9[]1;:Hc?B/7^KP)J[QV?a.(M^F:N4-b
E=<]abgNH[YDYLFK:Oc/?@#,/WdJEb[Oc&V?>5:FS:H.5GbC[Z5>2;;8a,FRd;-A
;:3)SJ1dHB.EQ\?EeJ92YOWNZ,70.0.=ZE=9XV/3N-\fc:Q24U[(NKU?/]a/(N4=
-(J2E7_@HGPG);:3,?I(4=)3c3</UQgK),6BRJ<M<(F?RUK8QR)[6HXI]V(I.5?e
MS,ZNeJ)K77F@X<7LPM^RE0#V](d=/\1ZG9d^;M+P_U_H.5I78>U8]3O?YbZ@-HP
X]D46(If)60@V891RFe@A<)XI&=;O#[14bB.\64;>.QQH?NJ8JPe9S,Z]AdVV&JX
4N&7,g^J96YN2.O;FC1WSO,DNHUUFGZ>>VU)^N#D)WF#.-NE(K6a^a6P[EN,_-S<
.61#WV65ZP8:4cATH74+2<<T,]&XgBDW5a=8-XN,:ZcCB>1?X/H].O:3>JJSXWL;
4IX9@M2AOE+Q:-BDMK0ST.S?^LAJ7(Q]&&X/_4A&Maa/f2a_Y/XQ0XY<e(4:@9SS
[AP#E,:b_F<f>S)-05&d77-^4;3;+VSJ3Gf+9a:_/^X_9,cBJB0A)6\;=H-GWZBE
,UIHNMF0JYEPU7:\T+fPg3-#F?+a5G30(-S+X+QCAb#+SLHK&.8SeKGGVZ).;^E@
P(B&=A_f.R2TPKWMD(ILS:NddSVa0]RHKc)TZ[IFX>)VFC7A8>:WV9HE/AO2LC0+
ZD@eB)eGEG[PM]BY52G7)d(&9TL3<:4gR1-8f_3E8@/:_JOS89cDB1-e;NW^/Raf
7_7L@?g\S+Kf[,eKLDB1)RI<g)>6Lg[.Of<3ScQ>J\1XbNW:N[c0^KbXCG^aY_\R
gaeP3:N\7:X:HgGAcZEJ,XV_-Td886_PKbVRGQ5JAcK4eX7gJ&=WJ?1a/=M,=1#/
B#IgCeFUJI#Ia^2?(1TH-:I/NH>#<-ZHU5.a1#Sbc2Z08TXR7RQ@9\64<V@[b+XQ
<8PdVESXNPX_;SZaB_/V<b/1Xfd[SXD[4NdTX0>b6[;7/69\NDN8^I(8Y\+YG2JU
5?8S+]#]BLdD:_ZSUDEX9aP5G)_1O3U6Y@DFW^5B\2;WKNLc6\<NdY8>Jf^T1XXR
LgKM-IO8NM\V1d<9GF/5=.Y)8HNB7O=c:^PJ[BHgFDd9R:R@RXH+#Y9RD9LB69&A
Q;(;_P)2@cQe8e6M3?D\<B4AbB7;b0=SN,(#8?<e]XBWF2=a)?JT#ZM026Z9NN(B
O/dCPQgA:I#MOI][B[.KG&QDd^O]b8OA=>LB8dfE=.F)X7RX31AF9(@B<?+09TW#
cC6)RR6NZ)R-;5^H@cV?H1\2H;aLCR[.]H-BL,A^LI7fe4FDGGKG2N[3c0c6#DKG
ccIVg3.QQ9@U8VfJ16OJdPSGL@f3WHFRC5:5,5:M?_1M,MJS;&XSJK;g(+>)?J,>
5]4S,E7W?AAJ<4]OKS:>V5PJ0W)0N@,6Z_F)BVc(Y+OGbKH?=0g4.17cB>aJ)/C0
9ZUYb8Jc+2))@@@S]^SQ)8/TEgSG]C5ZTg@[N6C0<\HPFH5EUVVU_gb0D1X/1-MJ
BY(//OCBS)AH?]>O:_1&gS1aCQ-PU=;KEZfWGfB<&](A3YU-SADB98@V-g/E7&Cd
-^4E?JNBd9aQ0H6:a/BAU-KMJ8,2S130XE)66bSWP2XF&I?S\)?5V#6cNg[X6,b6
I=b<NSRB_3?a^a-.,MeX>0W2a0X&-ePC)?e-:S30:Uc:<9#VGDNHdcR#>6;LD-de
/=KL-QIZ)PBW0=Q_g]5MS8[LRe/8_JEU;Le:FCFb/bb1D7[T=GYR4H;DW)T(.)dV
;9\]Kef_/5/(-7DUP9NaG<If:RR9&T/\1ce.M]6F&U<R>C2<-GRN&Cd,<LY)f#Ea
S^()UQ-(-ZG=6PLN:/A;EZ?I<B(MV3(T-:&.DbPJUPX7;c\ZKQ13L^]8AQNU<BA,
feRa5^;1JJKRRFeNJJROPAA7AD[MbfXF9,/0b(>U3f,M;BCea-0&X98F-0/N/U32
UfOMg8<a@MYG5aG;\,2Z5FX3]AOM@O1/6W2PD,@D+)JYW-HCK?H</M85YQaIO^_4
BH858>;L54PW_\IdJ@CG7I)PU#)+<L9c95:UDge,YIE<VF95Q3Ue.Q?\^QIA#fN:
AMPWGG&5D)3XaeUOJA8A[gDQWf7L/E2LN\7:6gcaCQU:B\0[KKcNH8b#616^WG:5
=>05+UcOE?EdEHf=JfVA1b]Ba)B+SeEDB[Z-HDgC]T2F6P&.5N_VVO#_R<+?-Q<)
LRT.[>)>).KQgWAKH4]AWOC]+c[;\HRP\EC&\K;NgN7IPg4<RQa)X&=1X&D4?8OK
\,M5RfL1BOY>a:/#9d0+BdLKJ,>Z[:0)7PZ/?b.JV>LXK>2ERXU-53a4+H;Pf;a>
?0D-^=E=CaK>:SEE2DB6X8f8H(a:Y]T/G:af#]TJ]T0PTTFSbU-JA0#Z\Q6E6K1?
/FQXXU.gE94J[\3MOI3K><9D[B7;W7L:6W918\OcF-(D@DbH29a.L\fF9M5:/-\I
S;P&5><,DC_H^?_4WW4,20KcHT>K[Cdf7dgH9b)LQ^(H\8,?[AH.,1Vc<RL6R<S>
aE71-#Q3SW[C_4C[[=?B9]ZIAE\_ZJJV+/@S--d</>_;L0X/[.DFUU7,S?@Y15O[
>M6_[dd3Z)=0^8E[#81UI19CVLZ+PGVdB/4V>@Z\>0=>:8)b3=>:eV&eLER19BGD
>(^c\_H#HB;/#=;H>QWcZFEN8f724C,W3OL09UEXDdGH<L;IZ/H9A/D/>WC8R\cI
c,PUcX4HOJ_g@Q>&)5/#d<OE_(8MWM#NddG3gJVAaXXK[d=86S-&Y6++Vf?U5P<H
[N4fU-g&dU)9<::DW7)T,VS]eIC@WBC):A@Te-/g^E6c_S8,Q5@d>2)S>#=2&+81
HQgO6Q5)XV9@,BbdReMA9W9.dfUHb=MVFZ-3GMRVT.G3G>\)/@J8/-BSE+dGeGA7
3:J,A.cYa:BXbM_V=S_MccPPZNZBH43@2]Y7<G,HING:<1C4f:@0?8Cd9Jf/&-8K
+SVRDOH57VgfI^XEU@&6M,;:-,-G416#EX-+cfdK#5>19<SJL,JY+f[)P&M.POLS
9a-ERHLMI.2bTP--?RD+.=-M0KZb^EGN]UXN#eB>C@E7g(+#4YDa_G;9.X&92a24
#NF+d1eD#Lg&Sf#-b_68&Y\5>\gTN<=e5a+3/J]MZ^Vd?K>A#]2T10H\=acd09JP
+7UVDKF5BU)CBBZ[_S@.7@TaH\:33,f@G_^Q]&d:c/Vb_F[_HdY:H4JZOV;E=ZE;
-;Fc[23)0&TgdQH0[Z51,DdY7\&-ZU_GOB#1,.O@<@K4E[CTQS9?;fRGTW?e>\UF
Ad,/5EU((8JM9Y=[Mg:W;<WA.GM]\]:5aEW.TFD>1NI&_H5ZL,BC@=SdDJE\?PR[
SLT^G7&59EJ87IDZXD]^0#IE&.?&COAafWV#95^;F0X8HJ+Id(+fTfM)EPCNO0]N
c^5AcLBfWHDZLe[U?A2<gC_QaLcK0Z_ALAM@YCC7^5Z(fSRV]M^XQW1SOZ7YRg#X
3APU=KHZJ:=:_:89]U6:R@dNH2_2,JKb8=;2R(^6\\e/\-eQ6]++:2>VII(DJPPV
?6X4J,8;bFd=&]MK<g][2a3PAd2fT(9@K14H<I8-fg.cb]-;9S>DL^S@4-:N>8cK
4HK[NY<^f:&gYM1WJ8Pe<^#Vb_LUa9-PPe\7CC#/PCIK;G(C#(-MFU8IIQ?)HJL3
bERK9UMagIVaP.M=?21.Q>;P[S+G=]KOd_WYO8I94XNLZEg;&8W(/Ra(:DR?;fY1
9e=VRX4g?G634d<E]c.[BLc2Q@F5N]/Cb.?#gdU\5T:N:dH;\Q9Nc0.=CQfHRWaW
@VdG7?>K/VaW[\C1@.8GN?ABX&Ma5X^NOR6#525CTT4ZIYVA0NZEE7VUDL8D>8S.
HL6dR;7GFD9J;RJP4\<[1&>&-CWg5g=EZ(4bG6:0KGQTc/GC#<Bc/5WYGbg9e/>E
N3(+EUTM&[<H]?+J_dJ>gd)5bf<[@AG/C4HWJ2?ZP-.L+1e#:(I.HL.S1N+[]@MG
@Q^5e+9DdPgHWaQFJ#[;\LD58N0A_7^8BfH6dL7A(YaLC7+YGReBgNOd>O34.-C]
I]gSKd#=F5:L906CQCK/:D9dWY82EMC@INg)^>48C[.92]aOAgGSJ):VUP2+HA,+
XHVdUNaI.,Y&UZ=>Ha2571dN.0fM&P?7HB:BM-/4eG0.91WQ]<f\XEc,#9+Z+6P;
:GeaE;A^]7D^<706ISS3)\UM<d:HdX<]@9cG^)?1+YLfEbB1gc>?g:29TGg91[H#
4e[&:=Z]X)X<;&a:KNX24]?=6N96T6=+QH.IF]1Hb;F1)dV82:P_,D8GeaLR+W8g
;&PV/1BX(1DA[F3>YSO;T+XXLfV0H-2MX)I]Wb=7-6+)SXG58RM^?3):<JbB#KMQ
ZHd/[8[,e=\^SRCed<18D@1DXE6E.]]fO4OG5SBaF-2RF4I4XTbO&8#6,DSWNccV
]SNbN/Y\S0:@.;J#7VTLQ-9VZI5^UF;I),A6PE+?)d>]/Qb[OXb<BbdWI?:)OJbH
f)\G3IeVRGS:7]3=;8M4Q9X:_b?I-cfdJ5I[Q95b_b\b:EcJ60SU\\GS)1TOY6Bf
2_IKR>O^WN_+UMAH,gU8#1AAO8Hc,AU5dGcJ]f&PERRVX47]A5WDeEGI7/CJRD1^
MC47D2O2KbAg:CB@8eAME#K@9/BBgAT6SM+5BKA>N<>ge3#060L,8_?8\gRCJgN3
;8b<7K.I7b[f9Y?G[US]_d<;J+&;TF6QVH8PObFb^O6#Tb.gJ4R5CZf_)5e4[b3\
8-0c)G?L]\B]f9^<H21RW&+8NMXQA()H=bVKaB16P(e^?K-237[]B+f7[61\C-J-
3X_55O_UX#P^).Z8g&^U+WGA#9=TgLBCE(E?]cV)P[3dIQ8Y^.b+_IZfHTE;L8bU
7QENBS1J>^;0eC)ag\,&,YbY2\gOcSZ:ZUY\^2/4Va.SBbJ^SQ(C\0;CNeca0S^6
>3J+:D)50X(QfN--;\\cL.1VP@PU?b@Qc7N9CR:eD>]8+IHPb,;@#Q5b+)0J_a:Y
AU,SLLR>a^HI.2Vd]/V[9#1^&46FeM,&.@OZH>.LAO@f&>7OF2,=M0)f;1cPQ8>1
&9P#bc>B=M>,<?\fOJ=PC]DIaGe:_-[@-EeT3CgQ,/e>-P8=_R=\MTV/F+#_^>HC
FOL(,CZ+,-U\a@SN)SGWO36-&;W_XWcN@/S[B#LOT-[KRVM[94&fTdK)BCXBe^VN
^-3?KDbR2)AE+P(f#T31W_4\=0W^W[CTfUCK#8Nd7\G-UZE2.M>GRC^IE=>X@?8A
9-39)58[R6c0X>U-.bUTA8Z.G^<JeBAQ_eO_[&(+^=:4KNT#FFNZ1bAG-LfY>W0]
611=#dU/5I-Kg^7Y,(ERC3ec33G3J]f+7BJLW_Rg-F^C=?W@@R1K9Z>NQJ5Ff;eG
;M+T6MaO>NY/Jf<1#^WS,TX@]^bH&\-?@?=XV\4E4+-AV-TH&)9&<-:dH3JR,ZTC
^NY&_B5NeD7H<OA6>75(4\I3PV\RTMC9[R\WQdYeOZBKf5J0T\60)Yd,OaSJD9ND
4c.F@cQ(9G;9/14)Gd#-23KQ-S@:BZ/.@T4^:)^4VI<-J5W;BJEFJ4(-=2LUY3-5
<cc^)N>ZF)_RcBXJRc.J3Sf?F7/OK+JX\_F[C;(69<;AT(6,&FGL,+IQ\3(>K1F&
-b[S\?FcEDCZ,85<AgS\g60R(?_:YdaY<CZ._56E[eOH>[&<L+:3dEDF4=T=dI7(
D2C)dD-^P8PCZ&aQB1\DVGKYM[+(CIKOCYK/(I,71BT1+4e\Ta1>>S_4Fg7:4WTU
PFY8GLIO2\XP-[K?.?8[XRA@-J7A?(#QGgcO&#gTR^?>@N#Z.E.+,NX8YcWN1cI#
bP[643-V-HIH0gKcB-6Z[)+,(g<e^?G8=+>E?CTPPM/1.R3)c@ZV7I<,>Hg0,WZE
GgYdI32X<6=;7N@G2B()C;]/=[3U0]Z3;DbJ3+U)e?\;XD-A(J+5NB>aEYXXC(;,
da=HH:#++H;638HI^I6TENOI@eb&OcEQ=a7=g5,G6d,Ya0Z.78/LI8<3DSEUISUc
A[8[:A@02,T)0YZ(Ue=bXCdG;@+XfN#g)RU(R6+W:/)SL[QOG[A1^F;G2UTGf-4V
;YJ5/F=2Y1[V\55&Y@D6MQV>?V5)ZLDd9EF1I\e8=1)e+8LgM,6V7)[_3faXeEFN
Rf\d0O,10<P/8HBW;WZT?&C3Rg0,PJSE2F8FMf(I3)Kd2S5AFK/#_OGHUPObOf@-
g+<QY\L\R.MVRWCV1AA@d&+ffJK);)RGL(N2X@1WDb^F8KM)5LfF<SW+AQ@eVWSP
7Y9]T]8WQU8BJK@\5&8O4YCJE7;/+>H4#WR;W#P>+dUd1VHdLcZa-7^G?\CdHXS_
,Qe.>23J_.cX17WG\:3HL=Y#,3P@3/F#JN0J@=M(:,&7=;LE9T^)CGN/YXA)gZ4Q
HNMNg6LDa-NWeL31X50]dRbM>Y70;)9D_gGFZcQ\;CRJ@F^TABLEE\S_BAK:cI:K
,9OWZ^fH29Y+\:cT-JefCU3)[>g:>,E)J0JW=)-f<I:;ZLF66HB47>F+K0H4OSG+
?8ZAK//@A13@TR1O4]4M4#/N_ac)=83>PeJ^H.4[+Z2&0#fO-0G.8M>JADH7c=_D
d5O9+c=Q&@2/^)60^X-(.[YG,MWaHN9VD=LDJQcX?ZW6L6Z[5U^[GNO-H,F)_UH>
4+9&a^8=D[cDHY(Q:^]c[\[eg).-^Zbc#cC;A]O..9F2@0J;Z_3eKRM2S3E^e@W=
30L?03U@WFW26AZNKaQ8d>+YYM)WS6XU7U>MK3FbCf:g#FSV&1e2SXGBM8KX,-?N
K/V:gSc[PBd,dQ+c(IOceZ]6#^U0I?7\FZgZ>50-0?1I5N(a)A=]8eJb-HV);?(K
]UZSW0=UQ7DEI7KA1LSVQZZ8gJ6R=K,258Dd:H,KQLMe5N?XA42HL]X2fD>gg4^B
;.C9()gUQ]a/J65TH.1Q41ZM=MBe#3-M:B/PWGFJ8Q5C4EU#3eM.@C^N/#.MaN<d
/<g#5_>AXd4[\Kg#&L:2(b1PRYeRKaf&c7^Y7c[F<X@&[-Ga,6F^@fM-48F>50(/
9=QUI)bQFUPWL\S-L([7J(3Eg]@I>DR>MTB93B<c3J2U7?<W0?V\T9E[bO_D_+]R
=7_MEX#T_@CV)MC\GELIUTb8b5df8U&M9>X79aV1YO@LQY<NeT+GbHF\LQ54SAJV
b._+?<N[AWaZ.]Q(b(.HXX3/c&5GM<JG];\KYZ-f9A8XYLfMgQ=L21G?=3F#6f0G
PBND3]<1Dg,[2U-O.[MFeGRQSH/eM3_P;6C=E[UVYN&NQK[=eU;_XTRH&]/N_Y32
c3d7H;QA9)(HMaJ>gW1HbPLAKJJ]&NHHbYaa5@RNL^D]XX+UNS9b:1G?1S#_(d2L
K25Y:FXEK#GGf&;BIe1gANV4U<G7FT7H7_KS7]^PG3AEM[bP=d.5f:Uc6M8;X/eB
N#4JF=(NH,#6,F8)]L&1P7.OY[V-e.Y=/DedQ77@Q6fVM_7f60fJ;10S_B>627f<
TIfESbgD-;LH?]fIA&NI6#4,U76[dOG0?#81d\A2(KPWNP;S=#3.H/[H#,?<1(_U
C<TfTgKBcE@+V]=LXX9Yb95R>LF;LRCQ6IV5#S3MN;AXW6SO^Ga^b>&-=N#0CV:?
L<_<f:+Y^/\(OJJd)Ie^G98bML?f:+C?F<;#30XQF:&^NY<MU9.Fe@Hdd6TeL[[R
BUAH1)_f9_>=f38#^[^bKA6Ugb#3]U=^0O>XNS/a_@LNQWN91]VXG(J\0U]_ZDG.
1<Y&H89<]:aM)/=dVA(4UB-6XcX#P\#E4@Z2+D>RN&<]WdV6cb.BDfBZWGUa/ZQ2
)38UOgJ0DR+SN3MP2R/#R4L-EbdSVeXcIeB0)5Yed4?KNa(Gea-RVHROgd[.f5=M
;IB2]]cV&Xf@Yb>E:a@\3H12\XU2OI\D[V[9eM>^,;A_&3XU>X0a+<QVbR#GT\.)
6U=c#^8\6[4IQ>Ve=I@0Bg@[be]SeG1FZ@06a?A,=[_JR1NX:>fb3]+SQE+[e<EA
cK+@gRTQ.6GX2AT:#5+GW]eYJ[G046BbXCc0OXa=N(-Ta3bN>P2dEC(S,[,]1_C+
(+]aT->)=?VO<0)J&b8J2X>T#:<Wdd,M3R=e0#DZ\8<H+\Mbb&Le<4\4f7=7Q9CK
5:0\F(.8F;3SWI0/IBM1PA@3G.c_c?F3T&:YPZ.g]cIC2+/U8Z0D7;_1U?U[Z5KP
L#-AGVgAW6#2_@cBJ8OJ5<=I;HR[/Q^8]QT.,;?@44^FG6.2C34;AV:+[\g-cL&A
//7g&[P)(P#+],X7fbWQF0C,eLN#Of\JH7d96b7N#Hee?GH+YR/RBFBI-TgX2a>C
K4_S[@7P,fa(M8U3<edXP5K[(>RD&POPU\2#@7L2cba0(<E2^(^D37T4gd7,R#[J
P@@beR8/&5P/JN&S0b+g4==c9L3&F@:#.^LdC[7S><1<Q@00V&L:08Eb/F6T50PA
RNOG<H3^?aUHXN:]P/DYN?Z)XX?F6Q=O7N+MTdYO78<aFc#=P1TC5FBMWS3#5WL-
O=;_U9#aX]fa#1Y]IC,aU-LU.WH(L,(Qc<a#7B7P8c(VJ>H:=S3_O1VX@NAF7b0_
egE,L#TD)TXb;>Ig7Fa(gYKU6B;M1NCG?5(FHHBW:@T+O?:J6&KV^J]N+=,?@=G5
gKB7b)FWCUZLW9.1JF[]4FSPLEf4#P5Kc+5Ie>#OX>Uf02?-Z+f#\#a@.CCd8#QA
Q])#::TK#-WDA51:;F[TfQ.N9N>6<A-)g&@DW>M_aJN>OeE?Ga(T4/H4#3,W1G[Q
0:<X1.(HdWMRJ^,J5#QP@>-=M;P;RFDL1:7-(J=ZPfP7YS8>.ND^aP/@:90ZKdLI
dQHH#OZ>gTCaLF,IaU:=FO/_?..3^4?-We-0KA+2:#.PI&@HMYD#ZXT51ZL:Q#f0
J1<f7bbA07C0Fg:aUQNAT#g(VEcd]W+1^\,>bF^c?^P<O1gT5c51IZ_Z_92>;9M7
eSY5I??]/4?=:&\<07-bCQ&JIZ=2^&e?A_^&]AIbdaXb++e9f)VI@1dE-;_e@G_f
R-bY]J8(R@_GR7=)B+_O5Kb8B^^dd][PLBdJD?@MNH.&cWgC3CW0Y]+P_^0SV)L]
XYa8(A(gVe?[8DP)+O@HE3>A@G#HP<&TVDB?(\A:M+>S_J_=29_4S\Mb75BSRA/e
E3;Cc?8>,59UR?@YG09_\6B#Y#BUDZ3VcVI/G]-Df6EWPG.7a4TGO(a@-D8>NX0I
J8,NI.]#2-_=TJ.1]SKUc1?SH0XgTR6=<_[d#N>D5CLSQ/?8H2M;8ZM2=g&68V5O
^M01J+7b@++UT?03\<+TM>X@;[D+&&^ZNQFJ4afQ1WGe?VW36UY7fIKTH<>(BOH&
G40Y@0RPGJ(Og-+(+\,<[bPBe]T=)K+7OS54^DRACde:N8227?6@B#^]NcSATe^\
Q5H_.b]FFBfC=41AEP+<H5A;M>Q(?f=I-DSNg-0a>E2e<WH0/[JZZF.geZ9WXM_:
,J.TY.TM0BU;3ID)KN?CVHdS&>(TO/JKc600Za;X9^FL--6N.cITe5][O91Y\I0;
.7?4]R&gQL]0bLO@LS8@,KcS6?X^a,M/V(85#&H(T\NY>e6+aUf&9;f7QHY7W9;a
&@Ne-YR=DU5X\Z^P4E.eM,T</LG&S[B(455A2^[C#6D-a/\D))80;Zf1P?5=?@-^
Z=eQC8DY+)Q3H[#M&;082G7M6JgPFHO5S/N&=^S=CH_#MZ<CBB7;gUU1KafFF?Cf
EXAg<]40G?>;;]V&4d9PER(33=-F[@>9ND<1,0A0F4)a/3U#Y870f?YPc08K./7f
K>N3,#>\)4B1C/4Q4Y6;KS^+8P-:3(OAME7+=)fKZ)<A_;bV5X4XQV0PQF81:QW:
)>g<?0J&8TEK8GOQIOCQQ&0IH3YfI8;5g@g5TI7+.I2#E06dUH3-R8F4f.>PSD&O
?^XScG4@7@.5J.AF/3277f:(\:28\DW#V0agTU,_J2(FV0P=01HY,1?PZPeCOOf5
G?8&85@\<W,YdYAR#B1JIQdcH7H0;Z.)+^Qe1D3A(GddGELORNbZQI9Z]28]X7bJ
#G]fDZdUB9/,TPOU(c2+O)S0>VRTW\CP2G[&4K;GP7&H83Qd_SK5:Bgb<DGF18PP
V_1>9F^S2OLf^dI[#c;H#b.C/)S[2Meg^;G69\F@MIOZTMT24f>/,B\2S/e=[EFd
U^:[8V04V2AL4@fZ^<\PF+HZYa(7#W==[GJ-GS1eCdgVI-81(XEN0fILAFaWaVSG
IT\VVbf3.J+<]3_6_NR.64Q<Kb#SSODTFA+LHb:9]LafSC[2bP@.<K\1([5c>Gf\
Xf^?M@]Vg\>W^8MR-,<@ggUSO&V/63:Pd;N@S8]39U;S]N+2M@TW.SNZJ,K]8/38
6NT4gI)e#8X2T\42,JO)8\[KEW(;M;1#U9:f(0>UU;L5+0R3_QVJ[[Z10T>M&G>g
:_#N2J>\G)4@6)]-9?PTC9KQ@,dTBNN>,+e<_<;+3>^dDfd(W.1/^4.daT=O-F6O
XQBaOIEc^?^(2@<^+^AD-/dQ0+MC1IXM5>V[,bE/aF]c;]DJEUdAg3,G8B=K,PX>
8MP:G,D-]@-;:&50T>Re)+e.J+c]&D6#Y4YS]g,dMH5^N]@3b+.^:XeF\\[?U2(V
9eDD4AV/40KePE4UGB<N[K?JO;g[d-55FSH9OcAagf[\LMGcf(447WN&0RL<TOU\
JT?UR#721Ybg>dd@UB7>>Fe(#OKMKD).305\ZQcRg1KgLH\#T?(^/O39Cf699KQE
4AcRQO@PfUQIWD0@c&&T2a]?LAIKQbYC7>3/Q^R;>I&B,\BH.A=a3#:;6CJCHVQ3
,P&8G[AcED#?B&J3Mc+&1ZM-UA\)P4Yg(5Be2[0a^Dc]#35,b6d_TXW\5b8@DP_9
H^5TZ/Od]/8HGY#9F_7?SF?[aa\b\Y[SL;Kf<(3::4Y#(F,93De1Fc_ZJD<VM6XB
I]P4W<W4L5F1&LVD(ES+,-WV+D4YOQ:>1cZ0BDFF=X9(cfUQJ^FUV[BDM<W&/]Z0
\WbWSSO5(__NHB>&X727g@.O=]W.gJ50Z8<9=gB,7=.79)QUW?9PY5TM+6EX]^J]
@f7M@NL.HR\MBPfS>OLATWe]:Z-5E)WIK+-7Z@RQ?M8J>,XJcN3(D3FER,gXOM]>
R4b(SV85O,OfXSP4S1>U8FT]HW12L/\<>RNDD/O]ZMXN]@P6U:XNKLD00gGR.\T_
H(9X-GA/JF2gEDU33V@V[XXR9R]KV+6B8)<GSf.9-U?^=V&KJ<-E^&Uf^&O]Q:BE
01eXPBdS<T2cIH/X^3/3=>AI5TVbX8KOD:\HI?R#LP3)a^&5+Lg&a@7Lb[UBBFd/
@FN:0>6HPPL1f#1O]FM7BGF^/EL9P[8I:RMA2FB-UA(_[;-DI<Q3>C;O0dc@)7cT
e\OGYSA3^YJfEG<3M92G+C<IOXY5\XB.T1M+#K92_FWWZTR<5.YD?H+:J>]Q263)
J<AL,(b2?3YA0LJ]-^H@2]-SUEYGNX[0ON\L6K)Tf5ULc5(0dTPCUV1GA:_&)029
+g,__G:g)>d\+Ue3.W#4VPI.9_&ZKSfUe33L<G1a:;:>gWMIC1M=:MCQ+C<P=aKF
QDWZ2O04>+;dO6,a=2.+J86[0(RP#;&KgXKJJU(Gfab<C08_8_Z0HNB\gf03cc:E
4V?94]3b4#CgZ9c3P6#\@4G1W+G#T;]S4&VU(U1##B2+JIZ\f,QP_V^/#9XL^Z#+
La@S01Sc13Z2]2<]^R1<Y3?/ScJ8=ONaAX\5d&EdCL:Xb2,Rcd;MR?3WAF/]?LdY
.Y?8=Z&)OQ9\@+3Z/CAe5==<=cPE?.b)]GfPcIa_Zc_GP6K,X,0H5R+.eW<c:\:G
-JK0-W]<c,CX?US97^PGc0N.[II;&1)NcHL)Q=@dK1IeIT\T&\)CR_E]#\:6?TZ6
b5cUJ?Q_/8&8^RH:^^beFbgV@T[aR3CDW9fZ<?#gG5GERD&3DJ+J5BK[C8_U=/N+
A20]Y\JI;cXKHX1Lg>X)fKA1L<E4c+X++&bAEOWH^DFH5eZCD=/6]NSL5Y<CG@.6
8;OD7VP?/ZAI_>^agSVWX,M2]dPV2WF<>I;Y]gf^KBZScRbB21B7<H:O06QgC7D:
b#W\Y)gIMOU;SS91JD[W20gORK:?]N/#BdPQ(V8E4&^(&/I0/KP-3FbS>-W]e/9N
2C>&)E:JTAO9?)g\-]W2&1Y)CaAY7-73<(5IIWO?0TYS6HRLe]^2WNWTILVP+g2^
Q#25PS4M_+[C2&V;dW?K+L7K:Z6?9;V-OSCK53;ILS,\&?c)3CUW^T9NMQbDZN[A
-JANb+cW+fa&&F<E=4-3aHN-BO@<Q#@;>2?a_=M7XT6)bJ0gV\)\bUSTW9c;HMB2
9IB<]4fL_^X7Z=HLKb#g>XH+>WdLP:2)3Cd47[/BEMc0LVfd94=^IC_\56_TP2FP
3G\GCO?d,@NYc6+Meb(NdgDV[+NP;5=B/;<d+.>ODWa6:?/2P,=5-TbW^VB?0-WP
[]Y.X1>c&U?>3<LY3Ad9G#Ib//>1W.@&+2eK:NKEZ&N^ZKO8aR(K2ScF9/GD1]AM
0b@-F2YQ^AeWZH9DQ/G>ZK9)J-PQN-APJ=0b:_:WW35F>X2_b]H:WHAVXdC>Xf6f
X9gXOJ:JR85L6XIF\MY-P7(/J2W)#&5Le33>Z:;bY4Lab])HaEcIA+L->+-,8<Y1
D(Vc]@-X7/e6A&O1N6AMIN2A+7(cEX\>YQD8B-C>H<OYHLN-67QM7d?;=U2KJAdc
\X1YTK;=<JHdgHRY^7d;L)5V:XYL@3+2;E\:c=0NH1RQ4a-HeA/LZDE>BUb&b<[G
aS#Z:gc6Z;T=XQG5eL;U;@_UZT1N\2(9#\Ag(a0L9>J4dgBgYOJ?#0b/MHQeO9Ef
.gec#S+BP@b\<84aNbDS[eEeG\B2Y;Vbf6ROcG?5H#>EONOAL-=,2\4?M<F..+22
WAGc5?\E2Ne\-D611(I8=LIJ^9UHC=?A\;)[A-MP,1[b,PdEb5+NHD_PeHFJ3Zd4
7D.PLW@?\/V(fQ3;g1(0g2Z#SN42;JEc9TA,b<#]?L^^W<b1XV\,JP_,JC-OPc51
d+>+94c2ff&T3ccaI(5LUeb/\HHAKPBMM8=9TX.)U\7+1L@H+1,(a]B51@6RgK82
N+21/.cDL#6W;B@^gI7V=1/DUBG>F_^a-eS^^:?_G5bV;Q-T.+ZH9)S4)NV:];K,
=[#e_@X=5TV=Gc,2g^E?1:+[_UYDE1?]HC>ITg42g(=_WZGH9[GY:0S<ZT?E7Ag?
]G,V2dZ@>7\0MH?(BbZU7aT.TMPeG_d8VRbT3-cFHFbIc)2.bFKX//3?:Z-]gS,Z
XgYA8KSK\HGdCH_UZ6ZM9c=,19[:FgJE/M6:b:CNYW\].KBUdg\c?Jc8PXF8aP-^
I3O+?N0@FNUIcGN(H79SgERf,WRRg#?&I]EaD^6g45f5Fd)17;XD5@J1QLBPT6b)
bK?26Ja-R+^ZU.MF,8d#\[\bUGUPJf;Q]]_2#3NG^36MO6VNKCVMg4\V\O?;c>6&
Y<.;B-.[X8d.XPCZVe>^]E>?b=V8#0Vcdg2LMZ4<#Qf6ZHC1<@5^<I9E])eL8,.:
Q(4TgRcD61<ZBWgc,-UgJ9/E6X<cLT62[M4bO=eM(A,=<CfAJCU>e)Ne1^IP)UAd
>Y;G<HH&/?e(@D\U-UOK.GY)\Z]3M6fe>NA73E/AdF6?<9N2T)6#_K0U7@8>fd^V
/G9,[>;WC185]Lf:2.(0DO/LS5F1]O??W-Z-6T]#M=1Y9Se\PNP3<4Q>Y_:&D:&Y
YTV=89,Ce,SU,T><#MN8O<_P?2=M)XGOOB460W+]+>;E.FN1MbQgZCX&8:(3DFTG
28LRY,9[B-QG^+28O4F)bcUH)<[BB0UDO36<L.fWY^VYJW5.OY55&YA[N\VRXW28
KGZO6O,@CVIVdaVP4C/Z2KFf)639b9SC<N8@16,US1e#I8]T&&aMLZ)2Z=+&e+OR
T\OH)Bd&BK?>fL0U-D49G?V_-(,X]?\CQK+9cd+dM^5f2^018Q)SIZVQUWZaGC;7
CJ&3WI9AGZ4V)C/[A=?0Hd\Z^F.bICI@M^/C^O4/U/4?e#G3U#e\b4P,()Y(C-RZ
@1,Hg)#\LAbF#>+Ie__,LOYF5TUQS6G[&0]2+3)@ZbK2+YE+01C,<TO3Je1)(-D/
MB3&-)cZaH_QQeP&7BI^R-EVa#WWFYM\bGTLQZQcY0aNfbK0+d@g)GG]4MA^3#dN
V@LZc&@)Sa0679da(9Q0KUD_334B(9ZSITAI/R)X)eLSV\+P6fF56?B>(aaT3:OA
Od)I7Y00ca3[^\Y1S<QMUFF@L\T2-_EcT-\DdOE+=MbNf<D3G&c5>\L1UUe44Ag&
=2-QBVJN#=<KL/4[Z<70fTaXN418=(-4b3IZ:,_<Y1PKLQKTL__e5]7)F=YW4M49
2DAK/1c?]&b(Y(+bE8?QLDOYcgWH&7P@UMPJP2QPONQ;NWUQLI1/f#&-a1<[cDef
9>Qd&):Y/[I@M:+fbX(5<#@2#7AIYGFS)I1Qc>e@93:Y2]D+C^bW#X;(BC&9?9+S
T_eDHAfLOD[K,RAd/B?a(WHHfJX+EIMaYGNXb\=--eBGUXcg2H.;gK03OSH[OI-U
_#&H0\+BP2,;8Q\95(AZ]Ja2NeA7S6HBN?MM/Y/ZL?3La^X]V:@04>D>d[4/?D1X
?bZ4d]DU#L^c7R]5d&K6)+:b8^GMcO_a.;gA3b<X3/gV&aDA46S5\=7aK?Q-)RCU
&T41\AV:d^L8TMG+VU.8QcOXO7+JdX_0I@=DHSFK&ScaPO5:a#]B>AT]L.9,c5#G
e/LZ+aN=?N8^gY?.1G<T?0dP.Ud2_3+f]Z5AIE8/dGaf65c1-Q(/^S,<A;4K(,OF
ZU2G9<^T&b#\.\N1aMb4).16QG[N)H08gdc3AQaQ[PQcMb<fcTEacc48KOfcM[2L
<9LJUF[/3<L6NMAHe@cD/3Q:^O5gZ>Y/;W@/JbFYSaN]S3@(C3RHM\f&K@cWW>^F
+#(:KRJ;76R3U1AOF6H\S&gF@Ac<;48.Q#32f\eXZD,L3D;W1_SLPHaWeCWW4J+;
.;eg)C7^,TW8d_ac#@44F&923ZP?GQdU9MW5]BLVG^K01#:2LJ2?<QO[,B#6_VSB
I7KA_[00\32Y^MK(P@K.PE#O;+BVN<G296=N>e#=fM5]eHZ;JWg:#40JW4-.N)aW
XV;HPWCE^-]\UWcAfZVC@.^g4OPB/.GU78):D(-D9_02]XG2<MQb?Zc^Wad3b;Qc
b#W5)QHg?4UVD<[J^/6=6.?D_N^Y4<B.Dc(@N)>8EI4LXK,?2XM,M=Q_4076gM;6
-e;O[EaU#F;LcgCc&Wc[[=cN<6-c@Ng.+\B50SLKP>9._c.6Df9cce1JcRNM#S5C
@WbC\?VDKa-8)Gd9[8;)+K3GH3#KO-=Z]BW59[8V.0FUKSB)D[\f2\SLI5L?J5e7
C/f^f9BfBB>30D.c7P&b.3U^>?H#JfReS,W;1BK@d4NbL:fPMSF\QgBe,FWVZdFC
LRfZ];T,G.:]>9YQb=8gMYTVGO<9Y3F>8=JFL70&OSF]A#),N&\b^CS.)Z>L8Ed+
DEd/P.&02RI((Z=#OG9BXS1MT_BY)c9^3_W/f/XAIg-bgCO)M)QRF@E#IWa?H@+H
F@T(Oc6O[0H\aD/-[UB<8fS[dc7DQ@/83QQ#DUa[ANg+WPaYGdb8&eC/OKNU@V8_
E/bP/;5B]A@WZ(YG3VC8e5GD[.18=A&4R\bJdZEJ3D4b2W2>MbPNcd#(CT5daZf+
=+EBT\9D?70@XY1F?3AC_ed3#9JgFQ;_;AL7_)@\:1g]>Ae-XM_dY?7:R<MJ[8@?
OQP[ZO2aP[AgGO)PFLK?:W)@&^14(1.DF:7d^].NfMZ&=[RCeC?.SNa80PQ5W#AK
92;;K<a:@cU-bR<\VegBG_-cdX>TJgD-Gcg61gGI\gGE.D<d]fT/)b-BC<00e:#)
I=<9/^&g)B0,Y<AX,0_^dgI5#A]K)E^g:-#d/[,ZJcOgR[K,FIe1RSGW<#J:<3?Z
B2BG__YKN6SK;+MeUQIfZ898Z\17UDfIEC9Z6];>AeM[SM)W;HEKBG)a/IS_gU_B
(ZK@9PJ5HbCVOEd/KT]bZ6_-W_[a@?@I3^U3aXc/fUU2CcESa3YfQI^T=^/[dTEF
S<8Ya]9.17B\DF1K.6>c,G:WM=DCN9L-bgfDZ/De9DH/,G)-8J,W1O0GAZT9aE>9
ePgL6\#GUbCF=,2@f3Aa-AVLZ28#N7bNJ/),S&E1I)R7Da8XPg80,PC?]CaC7c-E
=^AGaV\WMfA?XSd_aHQQfYXGTK7=K>4d8UT1PF_K4d:K-:D;:]Na2eeBFcD>bUH.
ba<B_eK-(GA(LM\X=RY-9UJ&;B?NNTT(1#2:<a=8@8?KX/bgEb\()<I/1@\KG[1>
3fI[9e5&^2^cF[<0V,.(E?(AT)VT8N/5VL^&)g/0D3J899+5_C;C(\>;QDQdd3gX
6U[ST@5fS\L#]??eRPCD:&ba=O-:gUALFI9/-P8>ML.S+:M[E-L1aB4L::3W.I(N
+ge1Q0Mc@OfCN:Z#58:OBfX^1f:93<DLD+g@c5_/9RTEDbPL.8<A.UI2D;aO^Z-a
?UEUKF#Y(Y[5CALFS6bDNH@7Nb2b.B0I[5Z^Sa&1J4&79(T^L8MDEX+7\?O8R5f(
.)(PPIWKNc2DI<@L=/+1[=Lf7:0D7L],1SIB^S.?K^=3=X4XDQ-A:<Xdc8ZOQc,@
3@,V:dg>7W;#@.E0b[Fa(7XUHWQQ36\9+2:dEKFQA6ZM,XMQEPf<1Ae]/S-LTZb-
MCgDB,Wc2BF((=8aVHRdc6L,9G36(^W@H);NJTRYXSXab]gYMN<2DT=.QL-CE8UK
3M<\YL/#_cBDX:#/Y#J[=#R]DEeY7a^eEIBgE]BZHKW3@#PO8;8(PKcI\LRQfZ;,
>J:,.JaQ<45NN2(N<DDUaHXc?8eeQQY=D9a7BfcR1P-HEHYRKDY^A:=1(8ZSd+^\
7f]&T](2_4D7?_+g+=]D?e]49V-9HKa=[:BDFF3U+K(Q;\(K5)NHaP-7H,O=K)Yc
O]LE31,6J_\:c]YIJB6L=ESdd+YXD_;,G-d,:fFE<^_De7^;KU4#WW]N]cd2d[==
@ID@e5Q70ZQ+,X47:B7bRfGRA&?RJ)A7_SM5459E]IAEY;fb(VS=5OQCYA&2U/].
PIM9b/Oab]2Dd0Kg+_F]:=WLXO\1=_(.C&,<Qd#Tb\@A6)4c=@[#fHU\IF+PTVB1
&I()R_W15Bg^eL8f,-cd<\OcDaKCN]2J5]<b-RRUWB53N2cW3CV[L)(9M/J(=A^/
8^53Ub()1QeegfN5egI5,G)A(d1)(g53DCK0+?,^KcEg^aP9&9CSUE9-&#R\7H>6
NQ,+U5Y3??-2+C68VE71MS6DQOKOeWMN>a])ZbUY=PG?af5+[-&@c>7MA@WM21&f
^Q=)RJ96Q2BRe#4JJ4+W\QC(C/IBaE.J9dCKAU&d+cgB>?YV+8H-)SFCIN](CCTP
DWTB_a=Z+F&ZQNC_L?#UOR,5NCZA4VS(3@Y@/&e5N>T\&g>&5<0MN64:-K7dH3A8
(RL<&&XZ=fB<c_U9d;X-C/OMXE8)L87]GC0AY83c5Q<0UT[KGK7#WXKH/:b7T^aZ
/Ga##4#K]P84O59dFL/1J1U4)dHMOXaB\3Q#8NJ98RX[27gdON?W]6^C@,?;,EZ2
f_OURec6[CU(<9MO8NE&_X5A5TXW:N9/Q20>H^;T(IP,VN)eMKDB#/MG\f]L(8V?
OROM#@,_<E_7;^2>/93;SVeXO0)\]PDBg7DFPAP3XO5?JBYbALV(@D;XR+5F[08>
YZ-.)M[KQNNFOCCM7^/#WSLVM0D.G4U0KX3LL7&T\\3W>0?=G__=FMc>d,[EI5&3
6^W_KC1R,eEBLKUgfc-VFIJ/:[-WJM,AVa.[3VZMf0YO(=L;-]R&F:++[=bL^[V6
O--=Sgc(KP#/TA2+Y[G]3Q<BgL4Kag8#.4RA\<e8)@Z\#d2Z.aJDW4=bGIWC>>.A
PT9TK6OJ,BX]BPAZIK7]LJ)4d#-4.8+_HO@B6,R.P-;;TYKRW/d;]/X.9]c->U8B
eUAN@HNFb^[gVNSL-AA8G=VGfcKZEcf=YNZ(Rd<]T_H<dJOg#>R1R[OY1P/RN2]_
b:cQFeG.7Ra^CI\?)Pc&1M(V0TP4\(,f,-Q-RA7dD=RfP,17811)d10RE&7O)g<7
-.\9gA]32SHe^RgSY79U8++#D0:RO\<^gX0gT_1ZCg,Y_F1RM.&G>dWX=BK2^CO6
,6(A\Q-^K=POK<aRQ:gQ^++=Ke-4N@e=0XLMQ..-^PMH>DWe?<W0+,I&DADdB/&N
4;?Uf47-:RdcF4BMV5G]Y]N0H<eY,KVV4c=^7D?Zec&,3]M9IC.S9UD>]C,<UCPJ
/O5f.\dN6HP4MLVY:;X)5GE^d?X&5=(:2Q;7H?(]Y38PR1VNH450TYG1B;?>27M4
P0O3TNePc<S:]dH=G.c@7HNZKT3>M:d2\MFH/6P/=>G^]Le#NW<I>9/6La&4-&X:
ZX+Kg7+18U;(IT,CYXOT6GXfGB>+][KMX#T6_B:d-AF9EFIY@US]IK&W15W]gJ.H
[SIN)5Oe5a3c6IcP(LaGM4^B2,E/;@1^gg/c[3XZf>3W9aO8-d#;:Tb#P1c)0:\W
A6,Fa&_.-PBbKP.2QHBY,I^g9O\N95KE_BH,=9KfGON>LD;6aHS0]c,A1I@-dYAI
?Y-WcSZA#EVA7OFdb_QF116D#LJ3.5TBa]9V)+0]E7HaOMB8-bFRV(1]>LFS:Q:S
S&T0aT+]1+R_^&[HgI@,.F9a]<^P\@NWF>8?B75K+S&RaRXUGP->JAB.B8>4Xd-;
\[OH&V.bV^:G#?FPb-G?0gO9O:JKDQ4Qda]F>R20S+U?4#:5_=HS?+:.UDRE-aD/
LI)U=4C.3<\X;NeT=Ib>VbbGd-G,dW,2\XUb&K<^e4:P@[T&X<J@3eGC>A=?Kf,D
P+C/MGKK)1a>0KH0-UQ=2Eg-HP)1WX(6Q[Ff/3VJ]YD2[7I)(:Z>8E,H[O<Vc_E3
3Z<3<KRP?:F_O&bKePDGBJ_GS094A)I7)QMTW7<fM(Za:+R2;<-6^YM=,?\f(4>W
?.gMKSE8dU#>eZUE5YRA_S&YDCXV:X<&]2KP>PFOg1Z6<@I+NbCA.^5A(?dX\eKd
AB<HRG6A0^c-SI5P=@,/]L557TV/ER[gW+E#CQC)X8&JFafD2T26UWf\NL9>EA#_
+RS3R:HLL)96fP&(0=bG0TVTXD#+TPH3\TS8c57CF/bgSe6>.#fe,VV^9CcGSOa(
FGS=OWZeNGWaZGO36VfS\Tb4<4.]PH&A7EU+,(=C>/3QgJFZG\IIX)@IPUbJA;DE
>UgHaX;d1Q+Q7O-=AdHT-:64C^;gbL>1]b(8J1dA-=^?PEI<a<d_]cAQ(3@]=5_J
bf[E?CaKU#>Z_A8B)\)/Vc8([U)f,0)+:JX^0\EENXc3IbDT1-8-@,?A<)\JdYNF
X&>3M1P>>WS1\_DGMP\K<Da0DP44Z@_N(D#M^S@fcEUEYb::/ZRHW-gU;=QIA21Q
+Q6E)9dF0JV)^WUA.SEcCO;(]3.;K,JDa?PYZQ]?^OH/WM:(SIJB._1M:BUM9F,3
ALfTOMM^4#.>M#9+;Z41?N,>Q2,J(FMIBa3K=/\DbSQ45UM/YY3Gf@;#0WT8R_\?
F=6Z0)CIVfgE[/#D:[g]g:41+X8HgE]I;(#O,QMDIV^O>QZJCDK\+bA=6\NP91=R
,E.^;>+2FLdHfI(4@>d=U@QeAM/5LX9#JFNBeB7Q\GJ&cQ/fU(].Q<1,=gaBB/;Q
<]-17Ma8.LX].Z77@X:POP36.g,.fPI,;BT2SXP)MHEd>B-G_5-+.GQH(+b<GGa^
FM+44[OR:U]CEK;CO.HU;-)(eOcbO7gCCdWaS)ZcQH1Md>K&GH-,@1C#]^PJPb]I
X>?@.S8S)XMAC:OK4^:]db/D_A&H^PWR4L:Nd2D#c81ISQ0FRg-NacO9)3M),B)+
WOHN9PC0c.D,+P6XCYA-0PdAPJ\UWRGSE>&CRBZ@3d0Y/SS,-)E;HJQZW>K=?L^G
K,d+22VR<LN)QgL/X/4cP&(J)47U.d(Y#9JX.fCQgg9T2XD^\X.-G\9(3[10OD.g
:MI(W7/EDK.<;b6SL<[:/SE.1]Y,)3JO#HYU:XJ;)>5g=:,dT:)3ebQc#DQ9V>@W
&f7Y_.)f<L>+S+C]?)9FZX\WSDaUUT8ba0:+-ZL-49@#TdGV-^_eX3fd1_EeHgZ6
#EcFTL=/@P&B]G9f^[Z@#Y&8_G/RFG>Xb0g&7Y0=IGg0@0:g4C(?R=CP-G0ENL66
B&9B@eP6PCR5^3&?#+F,HPZ_2,7Z)5\EHbT+Y^S7B9gZAGO^J4<IO^&<L2Z6T>:<
CJTQF]>Q8gJb6F\fN@G.d-TO+.FH(Y[a&cT4d<g^&?SI,>@f:JSQHdSB&U@,AdQ9
I,#&7e(4Z3D><(edC3L&T;(f2@5faU1c<Jg[E&M7<(I?8]:KG0-D0LWU5=MQ^29e
ZLR4PgF9>M0..N&/fc.CX:[FPAeD+DB7AIg;fY-<0.G>0_>8OKPXKEe8CY)UPT_.
EZFD:b5Hf,aG)?^@^:P/V>YM6a?A)L3?:5>EcX.3bR&IBK[gN5fVPC#B9H1a9DZ?
8&T16c6>:870T8PaCA3#bC>?B]S-+^NJK.37f?LUBdM)J_[>A4VdccWI:Z9PaOf]
:/>JE_0Vc,gbM+fA)_A,G<_\E.63b58(6U?(=[f.faAKb4&f/4?_-?=<<+<YS>+,
_SFJHRJT:A=3a:B3?YPaL5Pg#L,=VVda&#[P&A<c)]\)E<@-I?@\8(6>(U^,-a7B
W-&P:S>A?DI63IPG3;D-9HHV_)/9V>&&>IQ]a.eeDP0O90b:M)/=BgU\eG&+@_=]
e\,=6-feME.5XGA7](5HN49C_:>L>QX][AcK5(?X9XEZL/SG=-)4dC<]FQ:M;>SY
/0)aH+?XE\#S-3Jg3\A-&RXEY.+d+.]>DgXJaGbeAL__\f;[,5eBW@Bb=eDDfRVS
_SB)N;R(MEe>840VOYWBL6HHP?\>=ceP8V25eK&:Ld=eN[(4=RNeXMCN#7G,fX2>
/::B05)X35[C9NL__F8=GWWU)3G,[gT[+WUg/e7Q_]SP9VgEI)/_Ye7PDbIcId/a
0R@3E5LOdcSME3=09ef>OTAMKG3=@M\^@QgAGaUCR\5eU?)f^<H;0H0C=N_X)Z=e
#/^C^f4e71Uc/<E(W,SgS<eR7.#:2D#)=-(73#]fP]2MRQGe2&83PD5WHGNZ2=#T
;@/V#-aee&eNA#W0R=P&?3VF9M.bbDTe66f+#c#5<MVQ]YY(;SB01A7fGP9HIEfM
[6Y^N3SFES#C//>-a=A/BOM&;[_8/W)9aF2TbHHJ&&CL<UH3S.(G4e&G1JXE=3-D
WTf4^ROKPfXSTVRe7N6K7RO7^+HIFIQ/+]?/9G<O2-KZTX17^[c.0]a=0YT&64OC
H.(R,LB9@:>A50KN-6IV&Q^;6KP57Zf<9;K^@fM/O@7IHGW^:W;^2d47+FGTY+G<
/Pg+6SVP8>a8+WY>6VUa\X(G=gW/I>=/M8\f4g8]?4Of8)@Q0-eK/+]]M3&3@51g
WL1=aQA_M;PF\@gXM,>NVZ/:\2-;2P:?]QL.+51&>GC?2e[D109E2f[-T:ON(bE<
7ZJUPX@cS1815dV\E,+]ObO=^^IUb^dKFREY7LM15F&=J=)02-bH\&ZCg&3fg,1D
0QLG9Y)PHSU.2HX,M.6XLL4TaI&;B@Y[=F#-3M5ZcK58)Q>FU7JUNTCUAa;T6Qe#
99@98CK23b/#MbV]S4DD37c4D9>=8-;/#\E^T</ROP>caX4fca]:A&5JE6_UPS5G
^eW^0^d+Z&#Dc?;@R=M423;.]O7T<L.C8FF^3a+&?Z6U;_>g_#U0S?S[g@E-7=\M
U[/-3FD[)W7b76GJWV;1ff0]_EX9Y^XfDAE77CVaGK21TbF=^<8^#3_3Xg/?,S)D
&Gb[FFL-P[8G&dgX4,0@\DFD&&RCc&)bBH<,G-D5Z,4Me\DW&-]>GW:[>>\.b<cP
4dC8^QNZJ5YA_bYBa7O<8[?<O)/P&6W+FVXE_HcNbR>4X0AY#ZE]XP-\H[^CW?8Z
eb/U-]I+I?S?VBH>Yf?#]a2M=TCXZ,;fL>/&DS-gcZLR1LOE6(O:;a&N-M#@@6E-
(A),@._.L\UY=L9A=0S(^KMG;[Ieb<D.5#GCgH4:4LVP\M?(1C98C;-0V(#_D8.L
#U&^_;T>1@)R;E)LHbSHa4EP>dHgPfHc+J#X49(fD+c59P@90?XN>O-=H9IaKF,d
EU9)&OI?O><AUFUgCQ0#)cdV,+DFN]R=1-3\,1c)eD/8IX(bf?(\6FdBQa?,/RD;
:2JWT;[QO?TYRG0O^YbN8J=.82ZUd?CN1E<BW3OVK6I?ZHT#3Pg5WHA;@WeWebg2
VYM^REX.>),]W>-9C=R)-B1a@.Y-Kb?&95G9UeJ#VZ/fJLD9\9c<S.FS[X6Nc9(3
]TYO.W@S\PCXdZ&CW[BPVN@ATG?gAFY^WV,H4EVEV@H9g2/8gL<MM33)SF;dM3FL
M1ROUK=dENN+^@A3,?EBC2X(M0B7Ya-C@,N;G,H+BVcbECN@bS@aD8/e>MVH47]\
4&DFAP=J>@#<#b,<G[/6VaSda5IWXaR;9)_30fN1^Y.<-Ya#Xc+)#7[K>d\;dP[B
,^02XZeUER5FcRO[e20HcP.WXf:;/E#U1Oc6I;USDTXV^+U[8[YHUM,2gS:DO((2
\@A8):]7@.=Ka5X965LVURXZ9<4ag(2:0MY>=Ug25LCALJdI;\d0Y<S-S=HZ^U(V
XaA6SOI3P@YZEZVBDQUB3Y]-=&PDO-.I;g:G(1G-Me(d;f9IO&N\H-\NXYaDH[1/
OAT]X4#K[cW&E0T:F+-X&TF^:@abU7OTaf#;Z:W#e7>4N:C(I](A>R)P]73O&Jba
AC@G-@]Oeg;F_=_^^ZI8-(?XA)J_5A5SZ[+BG3,D(NeEO&AKc=0DZ1+57g1BXYPa
c,V4E.F5Cg;28VTW?-aBHL]cS+-(^MOLWOE=gAgH[GOR[QY8C\2I[#,C&LC)RK9g
Z]R[&6:,FBWZg?K980J[MTbK1]^VdeC)-0];-6]<#;C=g0?KT3W(9@8:)::DB#g#
X:CG\B1P^4>^6<HXb:IR3-b8=E6,f([R;J5N8Q9MV+1AT#U;A\cdUQ#Va@TSC#O_
:@>,IP?36Vf7IcQa?RS4SgET=8O.LBT+:K8[68M&:@UA-@S@QGbD4C8F1Egb:Y7I
^#YS.:+-(8=f2J+,7]KD9)LOU=AM6Kb@BV_3=1C5&#93\dC;7A1MbK(bSG;]41YI
/T3)A.[<2DWPWMSEeeY6+/@I^^(FV@cKKQE&R/(gTEEQ>cPG[-5Ra?.DF-I(,&A;
+GL/5_(:74>.<]#/TK68,KI/gPdbC.5(OM/)1W\+>IEUF@U^]Yc<3H(N-MI=W#1O
,QI0BD22]:EV\7SRdLfI7Q,E#FL[+fgL4:^<b64b\O#28Vg?XR8],]-8dBG^\f<C
<G5eD)0_9cefBbN]=0c<(2ePMBKC)]GXT9Z:c>fQf&(0GCEEV>DR@MI:@U;_ga3,
<9P_7WL5;/B##W7+SVU0eQ1J[>#=]MPS&#6EGJ/Z=INA0(?A5W1]]aMM+E^C<L7&
T8U#WZ\b\/L7gG8c8BJGV?>bC/CDVcYcD>B@cbNK6IE6D@-^2S,/1HL&9@_<IL.[
P8d)C]GaD,7^<c:K:8AIG/IfGb6?>X&,Z8EYga_f031S()WGI:dPAS7+XL#3d2CD
Ia@=B_FG3d7[-\]&=QfU4D25^T\^1EL;1G(K_fQ32^RUL+bYFMJ.MbA[<L1#^=U,
X6]]+CDgB_-YY2dJ_X9]QRgeH[\CB]Kd.G#gcgG4^.>^P_Wg6Y4:2(X78GSFJUe(
X5,+/<e<B:Y^@[>C\W1.5U=ZZ\7@8^04VUYNYAWa5[HM9Y=D+?(.aC<CAd(J&[=+
e..8WD3b_HOZ)g_>F:QH6^K9UeG158ccfR=6?fHa?:</X\f&(B+SM:.6C(3fW&0=
f;RKYKX;>1DK4IA@:YTC5JGQGLZfJaS4/9+8^L1F;fD1G&c+P^5T]WY@TH)T=&g5
eG@DV/;^UC<I=(\/;Kf,a&/<3D-aW&GX.M;H_SR9-2_>(BX^L>-Zbd3+RSaU_D&H
B)dVBY?=#BcN9c]a7F@Y9YI.I&Xc1<LKLOHRGF/Vf/dZS^EQcOER7Ec8^6M:X@e@
]M-[QS_VY^7S/N=SY+3=(INeK4K/&0K5Qa;@eNIHa/H+Cg4dNCWdX&LHBS>ZN,^3
efV_Q9<_?2<)SW]@O(QAbS#Dc]D3eOdBXdeK_a:=E\9aM#&aeM==\&S-<4+F&D\B
OQ.d2?QXgNM&S25M/#D1A:5#D6&IW+?4?U3ZV[VKCMg\\f^eO/IW2CN#5S<aL=L2
:_;Y];&5:CKY2-9gZ7.@QDI2L=;/03AG2H8d\^Ee_:aGS1O:OP[Y:IPEa?B)5:E5
AF8<4db,IC)C<O=WdM2_1E:cPFE]__6<Ue=@/>+.fKfAF\QOUf/T<-9R7M6TaRB_
1L.SYdA._W9Md0X&=>aQ6d3K2Df7)(0\/.J.(ZfA\e[eg?ZO[I3+J-/b92NTgGU0
ZY1Sg@CU4PN(Lbgb.bLL/@Q0M.7S4==.4&?FI3-^.?RZaTW,d/[B@Y,#]I]XDEX?
&W7fFZP:9J4J9ICPd7)09^]581A\eX)05C+=[A#U\#J9B;_Xg3<,?;ZCIH^Z?MZ=
<N-:J1DXOFdD;\R&.bf5D(R?\ZA,0/W[M4](2)@SSEa,V@NSL.^5/U@M3bcSW4>3
786+5C8Y6NMSa_OHZEN41_0?E9F7<VDA,X(^,GATQJ2ST-QdFE)RK03^\<0(;_-5
JCYV?Q/P-K8+I]/^d\T7CBY/-C8T/8;@[/g2O<E26WHVb#,be\C5N0J]_/)T<ad1
3OU#3C^MNW7G7_@).aSCRSNdaMET=^C=#G(<IO1_J,N^4WF[/YL34aE-1>>Mg;;M
e<XaZUc(4?.WMUNdL8Ee41()F8D9.eS(W;@SLVI2C(A&0F;]I>CP@906CB@e1aC<
PE5O81F]\41W(e-eP1=d@Y5e4SV1Efb_XYQ3OAL3+PABM<A1>B,fX4?#+D/3889V
P)I?@?587\.E@IQR&WL9X[]6\<Z?SS5<=(B[D&bd3E(/.G+37N@Yf]<>:#>.2]:K
7<&_&FVa2.4N2bV;K:g2VF\8COV\#U05K+0Mg0?]e:>-#bfX_TAaK[cKPWBc4SDe
W;[_PEYPWaW46\X:O8BSg-92=eO,URf\8aZX7&fKbdR+)+D4B[g5XTLGgZ9HK-P:
WN=IO;@A:KK4R,D])2fRNOCbF1JaJWEF6+C/W5Y5GgJ;c=+4U8QL;V[3BQED/L=4
\XdO_?;C<B8fJSE@(,_+29^De/&1:BBW010B^C1+CD/ZLBGK\;P\3[@[gEWZ.JFe
D@gdcM)&:LO\L8=:-Jc)?,6TMH#YF8<.G2VBGTU,#b9=3@;+3KdMQA5T8PZdg__1
C5c6,5,SK_aJ4PH@D+=X-A=Q^3a&X\>g)9JW(TAf^3#c)6^@D(.W>WbXL&MK+;TJ
E.4WEf/C+_?^,A@UN,W.Q1c5PDCIf(D&RSaIX,fJ[^:9ELZ.G2,SP,P];CgQB_0<
]0C09a<DLB=F/\NV34H\VMD3Td58\g-8S46@NY=(Z#5L.#gA+&?B#?^6G;PTR[I#
YQfGeUeP&4QU-I@@G(M)+aX4\4]&UYIf9c\UPTB-2BBQa[[3J3-TLZHY8UfE9Y6^
N__0,LI7Rg6V)R8N\_N)XV/@eeSF>J5TfOf&M<bV#5LPC0DDKe@IA;I1+X]JV#@-
MId_>AI:\8+35VCE9.BN+.U>&#X[X<3_8+c.0_bM(1AW:6-WeeD-B9_[R:1V/25D
U,e[ZJ?O5O]GDe3=D3M_8#0;S=547]cZ?;I.d&ZN6LQA\-D5CAaS1EG9EV=W5]6/
^UAV7Qe7K/cZcd+E8Z7CK\[2&)94[X>J8fZ3Y-_G,>d1Db9C??D,=/_0eEI=QY&+
gZ5:095+18Zg,&[:X-ZR@SP^=?AS>AcE<W&A1G\GDS<>S5X17[(V@Y5Ie?).F&-g
PWIHQXI^LMgFcX<1(-\HZD-R=-WU7;H(^I>/9.;deA2L]&O>^Q/a=-]FXD+DGJUP
LEU5J-#U>A&3-#I5+=Y+9@Ic)NCJe8A:.4dXQM>gcJ\&BeR96POe/I)ZGRHWY=Q8
&4DGHZE7WQ\_]MF2WdDeHA6CRL9PDO_L-HTRX;Z_:H&3bdIWJ;BER=5(O7fO5=60
^T3=7X_@]NWg/8a7>PMCbaTXN:Q]IM#3(#Q6d@D.Nc-6KZQY@RDMAWXaTCYKZJYc
D.WA/Y(,^[fMTa\?R@@ecBDgXI^6LG-f[2f[29DVR>=fJ2>b=KU?\_,P)K>DW7D^
g5K5?5>;>&fTWDFf+bS=gT3NRa2;QCe>+=e4Z,[M]MH7PY+b@E2a4e^:^U0f:^e_
I^6_:R].-/eQU?#a=Z:B1cSCJ5;WV,XK2UNL^[)E^(5N0]PCbC+6c.00ZP:D#b\Z
O?ZD?=K^C91-I;>6Vc4TW1HDN)]1cYW,,@H>-@I)Z(7&<:f_L0)ga&a(Ve+?<Mc(
.bE6NLL@NXZRPZ;3JHFXXgS+J5CCNaMTBV7bQY_=YHI0>:HD)+XP6^IYaI<]c\NO
VdBdWYW+P92(a10EX3X&+/,<72X<?2#47SR.M9]2Jabd<)g(aZG]4aG+VXW5c@41
aHOG9ZGOX)]Oe(E8?8\JN4@F;1M)fUbY\ZH.a+-3W\L]SQ.T.X/W8:VgE0aL4NA:
@[Z;RW?\3.]S_0/M48UQ<gYXSfF4geC53g#K#/aPH)^_&;T-4\-;HT,8>Y\O_G>O
gf_ZFB\)Be<@]7S3cFSOZRbDaMFV)<TL2X^ELBP-1QfAa-2?\Q<IM\U,<cD9AZM@
KP6LSX,[=3-L2S9b;)4C[7FH==?]1S3I^VXXfcc2H362;]3f6IP8M55aBCLG7T4G
J&b^X5:Y-2J8PDd=<W80YCPd<F(JbPG,/@YXRVeB\;<,UKZ3./d@ROWa^=#;AQBd
F@1CHY70.bRccCaY+SHXFEgLUW?#J.J9>7.VTKVe=g1[4Aa?Gb]&a7E>]J.9Z#7X
g-3A;#U>Rg=3d7-RZN#<LGQSEe,_><Ig@=gfN3@]-S7&C+)\2S](UdaUebBFV?fb
fbEGOgM4^>)QbY&3g1GQ67E.4D@g]@8-MM_,a/BcHNd6.+0Fb34UbTS]eO2H9\12
aYU3FbKfAN8Te:^NBXI=.a2)RD[2gd,Ug(]d(,ed&<&[_:#XV7O^ZAd(6@TJS=G4
gXGO.D,DAA5U(_0Q].1:Z=AadAR.5:?95g^3W^1XQ?A-1c7[(#Qf814I7a8B7V;H
^.F1^ZEbRMc,&@ZJ2.1Dc3F]^GK-^D:A&H]@a5(E:,CJ6ge[[)<f;D?:E7M=,:)W
TcU/];OKUOC\;a@<<18F5Rg4bK\/.TE>[48[RdDYQVb/(fR]aL\C1-YO+(UGRGUf
ZFUZ8-dBK_#(D(MWQLcMSRN3c4.5+[9=8BR3=cD\gHEW=F#]FBUK>D#W\E7dU-D.
,ZRO9ZM7<-D>JT;V145BJC8g_NMYNU/M=6-3DVP6&+VG4H5CHRZ;fT44Vc^?Gb&Q
N,\EQHO&9W2^\1&WYD;P<^QSRaOLC(Q8TYXdPU<11\@WR(OVRAB:O=cHAdONCF^[
</6;)UPIK31(\#M[-/:H(==c)M)AIQaS/Hf_?1.G2T>X[/d]_cgZ[;Kd[7TJ^I_4
VF4@ZWDW&V+CH@E,,2XA9Y8EB?)B^3@=\V55BV?\)eH#2c.]\]7-9GGZ,QXHQMF?
.?G3JIgCF8L:=&TV.ZAD+:Pe3_3.U_da],L6Z9/<R[O_1eX+Oc[C=PSgIf:679OK
,::I>H76Ga)];eW(/Ub5]-4b(;I>C\If.gQ[+_:K\XRN>]6;BHP[U\ZfaFHJIVZ=
gbb-N#H579gU/4^A^03a[:\-XZ/)LU/dHD,IBTW]]&.EM#=V3SW8GFV_c-Bb7eTH
<<U3[E\Z;4V\G1[b,PZE+#JA@g><@>;LCCD&QGL#^H?UFI[(]9ED_e\)Ab5ED\e8
3(>W+IKV[_FU3V853M)4#68HK,5=bDBb8C\ba3I4V7;]V?.G;Te\S+:A9LfVP&=)
2W[DA6]?Lc1]W139Y4^e2;#XCHFI>BR-#F1IYGUgW-8ZBAIfIfM]PNcg3:R=A#N+
eC&8a[.]T0TA?YdTRJ<QMe=,PcS=A6-5/OV6[IVOUP<4cMdCXCdJBI>D?DO?6+P,
#/,T+g#0FWa5b)=5?/_ZVQVG(ZJK1XG=,@V.-XZ=IVb\Fe<:Dd[O;cE24F(&bc^:
_/\)gPJ>4G;TI?H@Y0EL;S=TV4+U0Bfad_K\aZLJ4M;L\@?gN>Ic&/NHZ5@30=VU
@6Y7M24(TF#FR&ID-XFBBWc-?b04>EC1<FfQ(+HNQNfd:Ff4Y^L1F;ZX_B+)KA=P
a>(fFfAY_FLVLMa#6IK@CCdgd24OC73H+;f+]G[:6RAUg7W>+1-:_UW]bKZM8T2;
/27dJX0@JU-O7:>9=>_XTX:.I>cLU)fO/(X;DV>S4XKM_Hc8#\E@VE0GNF\XOU/6
[g=>fK_;89@X(#\C+[RRL9EFPR@N=LgAcB0K9(BP2)7K^bX+EQ184\(U@53<<;M2
J.bH3^6VP?=]GYDbaAOYSeeJU,,Y2NQ/WA0-d&eP;>WOY@-fc_[8M_>^fEYc)e9;
+<<d3?RSZOHIcNA.(bSN:E;QX^HD+e<>_#JXX88Y-;c([XcBGXD(UB+U[=I@>[5H
XC]b?b7VW38_9VR-bAEG/\K;Z?67,/ZJ/:@2Vd9ZX20>QaI3B(/d21-3T\</d2\>
Y(<Aa0XeD.G(0N]1K&Hb.[#JfOYG<(7I#D(9_D?AM:QfJ=X_M\c0/I3/B6fFCG2K
.))?ef61>f_QZ^^_6E0/M:/OVe/dB74JG9P)M0N\T2.:aQNF=8PFJcLSHb02U?Z\
1ZZU=/g@2U5P:(-7G>DR;8=\-YL+fR3:\aWU=4_KEK-JEP;CW+HcD5g0cVJB9H+7
VI7d:@_KQ@4-_7[Ygbe;:QEG6a27\,YW<GL0Aa7HBe6C0&TXA7RAB/g_N2N+LfOP
)QSC.WU?fZede<>ZGT(L4B>;gVW)7F+&/<01_SUbJ-K\YH4;(]\B,<C=e1A3Ne2P
LHYL7dZgWLYX9HDSg=V-#.@F09a-]PH^HFL4M.0Pc4H)W-Wa41>ZAK<Q;389FW^3
1,Zc7B((Z<1d;b^8NZGU1<^K67^\@g_/-<Vb@X_F(<Bg_A;FI.;Y83f]ACP6]V=6
F5)1cC[U<4&^<5KA[=GD:?&_df<X1<>[4PVJE/I]W[,4Z<+3M0>1gHA2Z_?=8E71
BE0=JQPaFa#]UJ^dgb6Y?N8EM,Z\(&_:2(YJgX&FOL2F-(GS^L16DL>KC8g63e4O
S6NBJ&AN^Q#-JXFK6HZ7YGJQcGKN0LKe+,W;M:LRC?._SM^H5SN49#_M=b[TeL4f
_EfMg1?O,N;@;fJ.C\0L]c;6Yb8gN1,_S2+W=g3fg0C(Ha(6RTPSDJ5=(>3/)>SG
3&[4>:#S+CdHVFF,]/2(GUC&=R,;d?RW0SKABG[TRCH7Q7A:TF)(>XE@:WNIgdbY
QJfg1FN2-^J#d=\MWMX@GU^U9?O]/+]67P4Sd3A/+Y6I_f]_\V6;Ta+E>F4^3^?F
2eCJ>,e3Zg3,9@&.+&@KWTOcc4@)-+]NS9<HbSF/K31XG,PT#XNN-@8,;d(N-W68
2ZOD(>]<b,I#4/aI>2=1VfQgQbM6-c99-gA:,JK8bc15934GD5.^4b:J#Sd4<fK.
4&;a7.,dJAS:ZZTBP@d8U=<g>(7/?F^g=<LBW+Z;[VSS.\g(?7H0-AVFdNX@#8cQ
PIfM3>)I\f6eN?UWA9S7K:)I8B;gT3M+VON+8bLSg[ES0dL.d<;1&D+S-6#(T]/B
gC0K][M[F@T,#RfU<3IgJ2U@AZ/dH,S/:HD[EC-X><,6XL4EP27Q-6N^8K(^VI/<
Y1KJ:KJ?He)1/7H,JQE4WB4CIOQRGO_I3OGSab\7=_JPKCWV0P-??.fR+F?[fT,^
-HcRGe+fM,:PPOc75[T@IIcPF/e8J75+YfE&/,MP:P)N?&aF9=E5O?EMV9^=TEYF
g(fQUY;)(;&@-S\VS3EX9@M6eOQ/W7:O02=C7ST29;SaTYP3A?8-bU,M2GOU\(7Y
2;(?^W(6U=-XB&_9,IaOL^(Af^8J-P[<]^c^9N/HD(OM?^D:Ce>b\QG\@e.2T7&I
A8B&^@X1BW&C1,S8g&17MG7?be\LCIK9U+J7YJ(4.,e5d+4(f<5?TNKP4<CKf067
\3:+2:#WII1/QCTMCb2f^/&6b4>,VE=P2O?XgL<?8OASB&=6K7NR&5;K>:HDFb.P
6?27)<-;BgNFYd[2.0gAHA#7KI_B/LMLM\f05TQCeG.OVOcf)5-<-dG5&B:YIT/H
#]^7A_=(M8BeEd-^cF>P<Bd7T/.A(:f1E;(<2^G<>G2b/.JLON-UF5b8..<FNTLQ
QCLGVFQ258EeECYNFV0BfXU,9+ZaT?2/_O5UNSUY;\#IOZ1:.+eMP<SEIXbM1PC/
O31S)XSNZP;,C#Pfb6:5-2H+TJIfE8b=I]g/:UF6^RE28@DWeEE8J<4]WcGQ8_RP
f_A.7;6EH6C;KD,Vbd@TF.V=13f0;/3^?\bWRZK;Qa\Yb@)Wc\M.KELKYPSeFaLZ
e#MT23][8)Y89Z736bH^S,6S9HbIZ&MSgJ8O+>L>&dQ7d]dIFMFVCJQaIO12QP(f
b_P(+C71fgNbY-1J#A?BL)+@X:-Agc37);1/U/H(-g/\-]L1IO3ATSB<c--T+#J9
JXZX-eQQIX^V78-GDc5DXWK=a-QJPWYY8d,+0fOX\#:@<2H0UMU3Q7<F)#FOg8G.
XG-Uf6##g=G96@R@ACO_:+2M+(6JD4\Z+Z-Z:SfVCbd-EX,N;942L:Y/PU2@+KaJ
\QXYYE^&.4OO\CK5?gWAPaT:/G),O0C8(JbJ^X5=^WMD:TDd;@8#_GP\U_(,]S9a
=L\[C1gCSF-7gT65KDAD+ZCRUQZg>5-_&2g,4=5=XS\&dGHPA]/J2/VBF8?OOaFN
P:W8/V(.\.5BOfV[4O]DE(d09EEC/H^W8g<NB,XI+f7BY.2-0g3K=<dLaD?EDcS:
Q+-5egTN(>e:4&KCf=9MQXLAZ\77K/I)_0?U(E3YfbJ#(P;/g-W5E8E5_:)DS)aY
G-00OT3A?XCJ?Ae05UALHf5)@M8WJ:M+]],UM<A.?8M>:)4K9TVI32SLcC.FC_27
OfX^gF5KN>+dW<Y<&3I]-()[,B:e()J->RdR0(A.P[Q=?JBXbB\Q6IeJLC:c,UWD
I&UaIY763@T7B6Y0ZA6aBO_6(<1.]RbJ)5Kb)AR)NHT)+ET=C1R22JZ?V/]1H&=+
KVS8XfPEI[;0K>b3#+)b<I>EP89PC,P8V)N4WedTA.8FXY7AO<dQ_YOB+gQ>eOKY
W9,<WEKCS@eBJAfg10A-JIQ/#</\Q&>[DJ7<KRAEH.ER<Sf;fM.42T0(3W7#:E3f
]UAU;4=/0)bG1WE-.Y#CAYc8b^S)&5ESH.&b#B]@5]BbQ19a8C=La.fgKV+4/(:g
:NVVfdV[>H-9a5+7#38GAL):\2#E0KL]@;EGFV&c25N1dC^[Z]80=DTfVE;W<^Zg
&)fYG_5S1Ig)FK1aVJN7>=5D?4Dd)>Y6/.Rb_:bOEDcJ;3EaHGeW.NDIa)VePC@L
0_fbKYEF1Q8d_@gN@0R+e4g4I=<I(>c,KI2G3BN].;7K[/9LU9Z87UMfRNI)JFcG
:aNK(V&E8RL,;e0@F\8a2R9KORTe(aX>0F0NAG-5gG)e_L)/9E_@,#(gMdH-5>V)
,cN^YY/GL)3#D<F][53BV49T/5:EeKe.C/LPJdd0(AN6?c5FHGO4M)]6WW[O?BYc
4GS/?7Wf+0D.)L6JXH1-9e8@[^Yd-[b1H(Vbc\;,T,E2dF8PG\XZNNWb_0Z;FR=1
]@,f-\J-L.ILLAK&0P@YB),a]/6bFd^;fCZN21/3M8[A?0X:RXG7e6G7K0EcFaV1
]ba?eKU(WaUECf-QNG)=P@+VB:W.N&#L39YW4HZL<W-355LJ=7VC3fJANULdDC>Y
dW+P,3U/UKfKT=8;2M+c0eYHRBY]VW0^&H7_E]a-B.E>a@IQGBS0T#_AS3KC:d]>
eNgNJ[Egb])?dRS/+\M@DW?>Pa=0P@(I[]L]WNZ;[)bfE#M7M\Y7RF>=,T++B2+(
YcX,QB0Y@\B,J?f]_0JG083.eGgLC.dIga_66140PG1QN<cEX<9L<1.ET<]PI(Pg
U()0M+af8U7>]<F^13)<&#9:Jc>>5=&I2N3c>VU++;7_\]GMH8<bZEU/bIRe7Y,;
;4301c=G?396_/J08G5F(-UX.fX1:1Kab>O):+-84_(e20S:H7F#6b62HWP7[?L>
>,1[Q\\11aa(U@ZE.3]F?I8Nd/=#YdKb.[>JHV;9X072gAIU)cEQVG6LC^D:c<\\
b@SM+<B1(EN]9d?1Z-gZG]7c:aJ<N7O[]ea#>4O)76AMa@2PJD;LYZgF@)Q]1J-=
beV-Jf#(@8D@6@;Q<5g>3N090&YE.A9F<dF[g=e[MFLZ6&R@&]#aMPQ:X//CLAW=
UZ]ERC=(.J8-fGf.5QC70/6f5_:^M3\_XHf\YP+UfAe]71^>0\JPWCS#2RY1L#M8
>aLLSWY3>,Y;:5F/>MKWUS:2-60+A+gg@DSJ(?BCfaf0TF&/F&d]F;8TV0e/:/K0
b^+,RNe,e1I8=<AG=Pfd:W^Q,&geR3)ON<b+,3JX[A&WXa0YSR6N5T=TYYY0)6IL
09b-O-<@YPfOQ+f6T2Y<efd2V[IV4\ORTKI91b9[7NaZUgc?d8;V]Vge^6^ac2V(
e6-D:B..LYc^,(bZ?X2S1a.\QeWY/bCe]BTWQ&f[7-F6AV:ffK(,DV2Z3#f<d2c1
Z6dL7(67):dUI+c)3[I@SYEQ6WNS)W>+L0S#4AX^Fa\55#9RF9T<8XWBML?)9O(g
J]7X8CR+EU/3Je3@S\U(cZ;]0R9N0KQ,-&5d^.JE<HSH7\1]Ce[\?A5X\)ZP]Ve-
cV]\MBFba+8b91352ecI2<baV_2^6(SPS^MF1MY]WCIUJ<APb_#HF#.\a4UV&c3J
&2W#eE[HG+&J3CY7G>./OAABKaPaVP2P=1S+5V8a83g9F^BN=,QY(+X327FYTI]b
XPI;(3#^T?B5:DX@bdg-dXAV97/&:C5Tc6=Z7bIE6fSbC)7V-\O&R#RHCd@?JW4F
3af;J:NZJN3F#/3<<Le[@_VIOb.8,?V36(8WKT-UO7JZ:=[D&0?Y,9X))]ga8fdd
M:gfQ4dX/cW,N?=&Q@\[0=9A5HBcD+:CH^MAF)b[OZYGZ&QLHX(2@?\=?a5XF0T^
.E+C-8ERbT=R_&>eaaOa(<Y8MI7<R==0I-aVC>]OGK;GQ;:H?19ID\]9,bA9.9YO
O_BLYXDHPLXaZ1QH^eEJU8a1-\5@,O/gQ36YT^=O;Kb^@S9J?<TZ(I/N^^)94GMD
[7(IW;SOa<<K6X-UL?54bYUQ\<+_J4J4a;HN2+OIU\.;]U\<SIY_XINQ;b^PGAE6
d[FG=bSEBb>PXBcI.X:4VJC6D6QIW1gO#I&4I^O7V=8GW4=bg>:6]5@ZdU,O?+g[
Ade>eg=eb;A3g]3\/A;G^DC\gNDH4QP?Df53-0-T+?I>d?Fb1\#W3^AL[9]J9(.=
,6/ZeR.6(Bg=DBH\ENR8#B:_^C<_:4-,A&P6#.^42E5aFIW=b@^16H0#E\]Z>d\9
A8eM>D]_2a@5dGB63AT6-:V8VAdV]0&;V=,,9VYY.b_D:?1/[4JZVL.d,:-bP?=[
2ED&;/R>\/F24UJegNEU:I?R:e\UA,NOQ_A/N-#KUYBNPUce_aUe&)e60P#[QR4e
A+(=I]P)VD8b,(6::<fZ;4+g4G+YF+GM5G+d+X9P9FAI>6Qe_P_3d\feC?8/_Q+F
^(<EBE?/+EfVL72VJ)]9EeCQ\gP.PP,1SN_\\L;+TVPT9\7Z/1[^0T:AMbQ.0b;g
^@(SQZWce#(V;<)X<>F89aL6SC3;QZ?1S4CWC;WVeDdL4[_MG7+@78U[.a.M+]+;
H0fZW4E.Bc3I+EDV6c8AIaMAOQD/H(&OF3X>M12?K._(]Y1Yc-FJPAd[ZHI+B>3-
IZA+X@C.IfE:>Y5Q>bafBU5NP+Q#^>O\LRU&\=?Y+[C[M4]Ia-Y&?LSP12CQ2Sc.
#?][(M<dYC^<.Q9P-EC>g[LC6Xd9J26_46dT7RQJTf@CMQB+7CXe#N3[IfFH:F6#
\FM\#\OWbBLU<,gU;T.1gR(<.U4C/c/0Q[N_OaU8S048YK_>B.JV=d1G+YU59-SE
C2&R,63]<M)0<E0V^>d@=cG<HJ/0<2Wba682@M0&2K,EK#e9KTDQ6^K-(=:QF+L=
=cTS:;[fSPBC.P/+PMegGT=\gI_)F7W/7Fd6^0NUSYS5=;R/?[RXc13/AUBT#KNX
aH=1YCQGBOV9;F?\<\&5)_J/>PS3:;R+VP92C@6SbSD.SZ++#;UHDG>MZ@F\R;N:
QV-/f;J-@Y<KM8/,DX:+GIQUb[@C1LS8Jc_<6b.D_gA)[E9B#5<_F\LZHKBI>3A8
Q:E=G_8<:C.L\JC2aBCQA:QVMUK=O&cfFAT6Y8NH+A-0CTD79WG9DV/?A-M[Mb)#
/Q7ZS].SYSbMB>1Y\a4=.,Ee_(3KM)(1^QdO-M/2.V)@39PY,SSR3b725<@6FX@Z
4F6d6c6gZE-YR\4>4<CFL_O68@N3BNA6(c;,OTH?)Y@>)g?7>X_ZNV#LEb7M=LSG
cfK#P<,^UCCBW7VP3063\f3^.d:\24&V,[Qb^EF\?]K^ASA,d<)(?#(-QKS-9.-6
_#[@c<-VSNAeAJ8I+F/7=(B=1#?Ae1/GR-M4eE>.M=.R8IF__G-g[?ae&SJKe,,G
d4<H/c&JKggAPC0WU+PW11XCQ+>[-TeQJB9f-;?2JXf-X6ZV_71@>f6:GY)1V;R7
<R-N(=7X16JF/CS4OL[T3/B:UL2/g+P7Z7IQ>/01KAF/:YfS=Hae[3J^55&Y->)S
=)^(3FIEc\U8LG[^3M]OGSC_=H?I.5XLN3&56)0HDe&7A&1KWe3#-A?U2bL?M61a
[eU5JbC^6N_@c\WK2<UAec)dEO<Rg2TE_,ZW,GbGe3ZDP_@e6EXMVd\_BD)=OFN(
2CG^N#375a>H0Y7SDP[R+/AE02#;AD2(5K:TAU.(Q,(b83\?L)\<O.(CQf[TIHPS
OZa+ZNQGB3F2:,3SNM\-;N\37G[98gG8.FT==:G++B##SbY2T[+5(Ke=Gd32OR)<
+b<);NH).\D34<CPE<BK>AIFW\D\g&K?<U+BC-CVCa.1X<1J#ggZ1ab(dTXg(F?d
fBEQ_3Z<SCK?Q@Rd=dEULe(0Z?c]^U^^BJ&IZ\GL5.EIX?c1<_(CR:D^TI5AU0TL
b@W9]8L5.6:WLYQCE=7QE0Z5CYWL5HE6OODG@\MS-_1Q?fL/+,4Z#L/OEVGN^X]A
eRU]8KP3A,V(-DM]Z8O^?P\Q:\dA&K9VOEE5YLT(@WYZ07:bb:UA3c1&AX[YNFJ6
ED3S8G?A<L(=26K=P5[3F>MDY,IfO9Rd&,8#),,QPU.TRS+-e(3,<_>OM)J]:F<9
4>.MZ-b[L]PDWR>Xd5<Wf2dC0OX;3,.2#^Y#9NUOK5Y5R,K,BMZ6F9,S@NeQ-8GU
Ue(@@[B,Ia4YK.HL]Q?_1eN>,1YU1))BN,9@WQ/2V(KN4GB)XS#ff)I-8[>5VKEH
D,?/L9U1CQN9=aMD3[;@W(ND1>(:5F>^IV<>-H->BO((a2#5W@,:WbCR1f1WE9UG
V^E+^LL5MK)?8c^XHOUfV7([@J]D&Y2Q_NJ7VN6QCD=-)+C;-6d[;,5CL#^DWXa0
)CVBXXY0D#;W];GC5GB[N<TEd\e?A+QYVF+F+>N1.+0?DA+HNJ3cb4PV(J#0_BOc
GB,-BL)QC.HMa,Y_#0^C.KB<V1WG8J_U(TbW5BM8V]H3E2&bcRIa.:\Qe36c58RA
-Tc1;X&V#T44,+H>/)1HUe9U_;Hg:SMW@RN#?KeZgP\2XPg9<c@0;?-e-MLB0D8F
NH;VNf^^VK\3(6+AF_);Z6MT6f7CfED@PLR=@/^=PS:.Q-PAUfX2.cG,00/8fC_?
0Gb/Q,S.1>_O[MbH(&S@TDS&5#LV08:NO.6T]R[g+S@/WQZ5AKA+fFUYg,37DBP5
&@@<#=>7(5O61A:VCD,[7XMfbA9U<7LIfG8cS\g[NNB=OV4PY3XGY4R+K\)4^TAL
:X[7cY):bMLe\<d7&&#5Igg7[@-EJ^Y6CSg.LN6&cb/#&5DMb.+dF]579FE(.6a0
L[R4Mb_K(cOg>J^5U17MTe]UAD>LLL8QO.AXf^g:g:2E08g7beOY2f?f>]H=[:\J
38\bZbPC5KC2UA<g3/J/>9DSCSR;_MMaSVfV@O127QB.^cYeZ<a6W8H5YT0/d[3V
W][<N=?)Hc7AXE3H6CaD?=0=d=1Q^L0E@?Z7a<e^W)6>U]ce+cY>)L,UCPD\(3Ed
06KF)9a^WZOMI3O;7aZ8[HO1d^DS+\<@_6edYJC._C@&C4O=f3[<@fXQ_M#b>/Wa
<.8Yc5S.7TN@M@#,1BWH@#Q-6H8#M/^;N]M=9[WP5B4>73L[\CBNR@6A>g+@ZNaP
Z9F+PbE9X5[80f=LRQ[EUO8eKP/95C(1D.04Z/9/,.)9dCV?W(EH]gNTU:5;OLcf
F,(,e9_(9RP@5F+f5ge+Z>T:RHf=aKgBCN6PECM?VgINT7))/NZWP>][.eOV9^.f
Y@.,8>NU7RS7GH0LeH:D)73SaFJ&-WFc(7F9(#5EX)a(T@cR9egV0N?/=30W+3:7
,=<B<--69<Z9JKP+O-:-H=)8()f>Ucf_JS-=7=R#-f8-=?LgODKW@2C[8E5Y5:c4
(GR>=_Z3H/RR+g3P#4]HV6-9QaU]R.7:(f/:X4C#J7O->aa.C(gRG2f[H7_gI(^S
(X\A4NFa6H8_J4SaB+PKWF95K>+#44C(;ZA/[MSOI[b1R7O]@Af38>WF_4dE5BD9
80?aO1]F[aV&YV0<>faGFUR39bf@>?MUZVJf[.L3NF?<;E2b^a23J<6\[CQ:-:_A
:R,dQ/3XV37Id1M-b#KCcB2:O\JSU,e79g_8GB^_(YSBVcQNRf7(=D;;](+;&&+J
FG4e-/L5a3#QG\I?ad;\9gCE6;6Cbee16<)3PAF1F>S:FSc04V]dG5dg^gUEV^J^
88b6E2+6U4E[c9N7ENH5M/+g.V&D(g@CTUeNF[0DM^,KL7ZX54R<T>-?G:W4FZPd
61Y1FWF@?4^Gd8#MYX5//QQ&#.QDUeMKb#0bFZ>4[aB-?K?\8WP1WBW[BL7_ZJ6H
3YF04UgXe&bOZgSO?:<gA;9@gUK9R@+(M3fdHSeDR^]#c5g9;LZ,LLEf10b.KdH&
;Z,Ka[B=83Z2]1ZRUU]7,(1R8gK5<XUJ<RLOabKDJ-70J_U@J4.c4@9c+&7O/4SV
3HBP+9.7,-b?cR&STfKfd/Yb9,(PbCfCdPCbQMa<RM3AW-g/T0M2\QS\67XM8,R#
e+U.18YROIXL4B_(:)b>5;3/O)GcS9D@.bWH&MYfK[Md<LHc(MX\GWP>5f@(;+bF
P:V+[c\Y0>VAU>.8_Yg?0JM(--IM^07:S.S?-_GF9Vc8-EK=P,K20aYGES(TRMOH
)e^_N_NdUV=.D(FZ2VTe(DCE(=FKU:f)6bNZ9<QOA?4I@(Og2>b.Fb-W3U7HE=MK
/:I-CGbPb(1+=GUUeM:b1dU5HR38ZMG=J</J/[b>]7KZG<K(G71Z]LC&D6\J5;H5
;.dFCTb#/d>1,XTG1H#e^f0#eU>K+[ZN9VCX8#XXS6c<C@<Sd?>P1)g^Y.:,e@Vg
+-EC0gS-YPW1c.\bW35>.PQI+Q).CNG8KOEF.,4V/\ga@I3a9>(Lgb3XHbO)0+:#
MPWg5Z+CZ0HAUGX15^f.AZ-2>-FPKg@[[;I3N&Xe7-R@&fRcM8ESFGC>3=3GZdLR
b_X2ea4M(AF.H5dg?&b?3b9gOFI^RL8L8e1:<;K#.g=6:YCb]&(-c]AVG-+63K^=
BAZ.<_3OG:LFQJ9cX6I)4VV&R/=FI<HB+5#dG97E3,?b^S;J3Z_>5ICENQ[Pd(BK
)6>^GQD2Z1Q/dK?UG7ZAK;f<9XBGb7/[/ESFP8.A]?I>a(^gFJX2A(BD^6DaE;4Q
PYPNJP1K[=H181LP#Q&ZO<ZF&BXPGg163f7#K:G-KCGPgZE9-E?Y;0IF;O<f89(G
+.9\I&DPD167B]IdL:-Jg3[/VR-)0/-82A[ae_J>1?DU)Q83?1T<##EXaPeEH>6@
S3\K)2(;2d[CcYDDAI(MT(O>\3Z:)78U&)P6#?H.#N];7U8?YBbH^)9WU6f/II^f
932@eG.\?bLNSW-P/_633Wg<PG#U;OMJ#,)?6XJTO^<L]S9TL-@Y[X4g3[Xg_b6c
S\)EbUC@Qb3SWS-:V:NL,@93cg35R1abO/P&Yd>7LU0_2gFb9=N.gXAe1>O/7U=2
NX)ZQYK1FPg]UX&SC+R3XG[f?G3B]?2M8X<^Gb3aEeBN>H<cLK#Y7,M85Y]XK=^f
#7=C&=UHdT,8(3BXUKP+L81-S:a/R40dTNcd[7&;gDPZDCU6M;?&Q=gb5c;K]8(D
GB2U-&HePMRPY5@36>+VRX35B;Z9][3_#a:X=MWG&]G3V/J?\/K&6XFTKSd.\)K_
#eP[\AfO:\RD@\.PP<9c>>?/Eb@[SHeHUWQ1@LGP)EA\=bV+]X\5S)+XJZ1EB+5?
d/+G?UV_:K9B-D?cD/91W;9Q(O6.),M]95H^1CEHONQ,WD[GV61DeQ[fOR?C(RUf
]bW+J-9(699(3Ic;4_6?7\K&F2>64W36c6N:XMN^++).S9PH,,?Na+MAfCB[(M#;
fXBd9EHG^_._8ZC7X/Y.LRL\Wf5L:AebbOOd\b\UMeccAY^A<[Y]G=9g:LX/G=Bb
;/&X&0KUS@fRJTXb=aCX7)S/T3TU,S#4VcON.F,&LLQ;]e7baUSa=[@(-3#YdN+1
e@?B4;1FO9Q5RT,L-]\3RUd>gFJ0J+]AFNXG)/g]KdOeB7;D65f^<5TBOaN.BCb?
G,NGJ>OI=)>^X(85U@Rf&WaO-g:VfNUa\#R;Lf8[0]-YZG-?bV&bLH,;K.&9P&c(
@)D\QOb.e/+G2Z3_;F&4;]d:TEP-@&</Z2)^>Q[K)8&I&=FX1H[T<g=OZ8a3UWeT
4CB(0@A8AJD/@&+V>TGcELF^Z#)aIMH_OIUALGaIP5?-Ea/03^eZ.P.bDE/3eg&=
+IMId[-R]Wf+6aCCG,>]JVJ0CPA7_MCMDCHV8=O[Q>MR2,@GI/9AMfA#OOSMJ52?
ISeC0&B\/]]K=+T4@^D8?UN@IgGPX\JL:4gN1b(7006W^]/MY5)V4O,LgE(a^17J
L5XaCJb@G1bW8f08c@.Jg.42Pa,589>KOP31]Mgd5=OUG6_g^-\TUKDSD]U0O&XG
LEcc:3\/-ZU6Mc[bB59>c9f4LXbIZ9K859XJ(FFb:eSDMML_g[4R/NY+6ILa\T/=
>a&U<C09PPR4[],.C(6G#Q;A:J3/=@XfQTg>X:Y(JNZW&@a8ac,XA>6QKV.U<,N5
=#;82)_BKM.,^UC?E^5JXca#d=OT?&RAL,D&/Vb;FR<#_(/@7;6OMbA#=b)H]RK^
L2OUDga=PZZ-He&V2BUSF08+(=4D9bN\J#&07dQHA8UBZ5TH7]F/(?@6c6Hd=06@
1,86LR8,f:X+PYf29-\^gg97V:(ET@Z-E>WGNeXA0[cUWGF(N0TI[B@L6Dc9.dgO
L;Gg8=1eLY5B,VP<>gA-HXXB;aW5^?-ZF-\]gHL@g2(T=?O4E1A=-D>0_HP<N&+Z
b.S-5EC/:A5UPPD(SCAV@KN)V(TaGS9;NWO<e+3>_W5DU#\B?&Xg9FW+U>,KBQDE
d_<,_40;ea00P^357e].c58[..TYA87)HXLMe7SB_-#):#O/14N54-U9ZCN5BZ/g
,0+a]MQXRfb3J4\;^)GOK_QHb-bAAOf)LFR;aIYbVD5RPdE\S>4>=(ID^=.7gDL+
XGCd>:=3#_@EHDd5FM&Y/7EW3:=3R)U&+V)Ze0,Dg[>+U0_KN#&aYEP?1(<#.UCC
P/^S\[&\eZX8B>.HYE&2R?bN,b8ME/L/M:d=DOE:fB5RDZH#;Z.]U(0<MDB;:;fF
1-H8)cGA<Y]bBAU+Kf?1?A[c3),gFY8SdH1W59M[\Ce@@>G=XHT3D/FI+fS>DMO]
)aBRDM+A>e=W1a_G#AT7\+V9g=\9f]]+/8M<&Ya/K52;S,J9,K<J,[W<_#OX35eK
7H?<1b2L;II)#K\2^@UQT@CWLFSe?>#G0#A\^:\9Z[:0-bY?I.b(+GHOX.8<@]34
BLAd.Rd?:HB<Zb[D[>[WX:J+H>TUW#.N#0<f_9B371;83WS4#d:#aZUUO<XQf+0K
JJ+Q[T0[.f5BBLD&X[HF&XK,Y[]DdS^M[/^Ye]TYK>[?.Gdc+(X[.@e8:#R];Ud;
bS?EOZO#?1]E.HTAgRg<d60:[5D810(T@DWd:NC/]K>a6b,6S-+[D:]&UWS)X)/f
a?_K;&.SB?^Y[Na+D^LMdUY571F+?[S/G@83-f.+59#UKL6MQ5HYI@;VI+E(K>)\
)N-fD0^@0M2E13<CTOZ^EK&WVT#,&+A)D6c0[BEW;?afU+1WSZ,T;IO5#G&,,CEb
Ld,>5+F]gXVZD^fC40+58F.^b4.UD+Ye)f0(OOYCE)90>(&Bg-;1eT\>d_4Q<+4^
M(57@^1Y;b3CR:19NI)8QS.(VPFbW&CbQ2GT1H5N@_=N&f+5P8POZO0[42e;e1S?
#@eZWff[UL-..]d&NZ8Q0UJgTBJa1L:^7/D-LbPX\7T<V<V+PdKb7NC7[A(08Uc?
&Y=B?PGH,bPX17;U<e6&\HV[O9YJda2(1=CC\34S7?SK]<@+O(^I/CRIfO2IQ9Cg
?,?Ne=36F9/L[_I:dES3_-M4G@SZeW&.NC\K.AdX1f.NJRJ\=Y6=QMcX1Zg2cC0a
fXJA84;GU=]@&PW#)2e14H/2d@#,\S0bJ_#(O;KJ4-FVV1#OEefbd,Nf9GVXB/@^
3M&U?9>B/L&+[Y-ZE:4UK-)+Y-SGUF[KGgUKAZUYVU-3:;g/LRPD03[EcIP8g1E9
c7@623B8QS=@<>P#G[4P0,c?J_[,>V,>,./E0KGTZIA#\-a>fZG52/G@&7b@G\MD
1CS85KB(af9AaG?#2Nd>f(D/eK]@TL8JR:NXY:8VLZQ=R^8fLV^;Yf?gPd?+dU&J
8;,21P(K\<)HD_DI9-XDI>[=CMLKMHVgLe,3FMO6X98G_-WY1-fcKT&D&8KQ,A>;
>=:\+X<?P0N]e0>.ZFdQ8V64X)33TE2JFVK;?=L4+U93fa@9E,779A;f/NU2C8>e
?R#IaA_3-Z71BOg>\U(g0;&&gV3&/AT0Fa6A0Ra-/H.&aJf?V=T7J0#P(M][(89I
_9dN=-&D6=3\,gI#@;deYK=Y@[KL>K#2D&ZdPAHJ<YX1\5E2>XH)4\)8^9)@C+6;
YUg48/IKf10##<JSUc,DdX(XTDO4K::VC)aC)gZDRCd#-RA//(Y.)C7gYJJaCO_W
G58@=16gEG10B0a=T^O_e(;;7aQE=Od]aY^)0]3;(]]G6<O0aE-B&F,c:+=F]WO&
aH/M7&VNP--AE]TRY2N6#=DSd[g59O_YZ@Eab,W6,=W.5LA:LE:REdF_(U>\HJ72
d#0-I\1>05.](Q.B9EX1@V.fbg#^-46CN-^-_3<YJ8bYd27eK@DcCd];?LK2R?_@
1\ddbGWfY]:)4C(<LN5#?eUbZ\S\Q/;S-T_([SU+A[\b)T;OKN48]@Re60I(G>FP
&O97?TG-),H_WT4E;4PXL4:,W.,V0U3:=83Fg#(G(L]1GQ-3eAdB1?O_JW>(?3b.
.<IU/<\g1GV;[_W;C#?EI?b]N-_c9T5M;AP6bT2@9NKedG]5=:NBWQ>HWX@7/K_Z
]SHHaJIP702c^e63+f9\1R];f-\/-EV4GT5ZBB.R:#L#>RC[;FfaJ_L:@SL,?@?.
^GA61e(<<@ZaZgbF#cOV;=TWX\>L3X1HD3,0\U#4QFU;a:eMS58DY:84C(Z;M6&D
cFP-;&[5)(GCeD)M#R+2O+VF:0_>_3;X.[<9G6a^M3,QP+=V&Vf,3/a3VLe5]eaB
_18f5T^g\bDMO_O#bf1:#UP)(V<[_>,@5[IVJ6J9N&Z55\QDg#X\)7+0F:&_?#L6
UOXPZ-JU,;FQUZ^CbT\,SF>9M[EFH(6(f+XW,VG9#03aXA,4cY=WIeJ^[\<b:C,S
6dO\A7<#?HdZ=d=2Z:gXg+b@5=5B+F90#SXOVXWN4Gf.8B;:#Id80WV1&VZ7P@P?
RD:19:e(ZQZ/9);>bJD[b4G(2?(@<-(g#][D8R@6(6@UP^cU2=Y2.WLB)+aD2<Kd
,XOc<ZW.^O7F:DZTGabB18^g?W=-?N\CJ\FQ</<(_g\I7C2L?FZcLC<M;#WNIbLF
.O-]84J[A>W[;f&1L6SNT_5H;DZ:f:\VaU>Mbe-X=[RMLc2bD\D.KZb\F>;SG3\\
/8-+_3UZ[ZH<&+]6[QVHHf-?V>@P/7=[2D)e:?3@WEC3;BK:?/(I(R2e;5&==-?C
Z9N1D<QB;[RIZE@<:Pb#.9IP)JK+W#+b72B)(-@LQW<1GMN?;a5fAADO0LH[ZbLC
R24V:[DP.1E_^g_Y?>O;20aB:.)g-&^-Sg:bX]2e+bE,b:_8ZTce]^^_BH>OBS2B
bUGQ2O3II0ZeWSU0bfg?7TTI@Z&:)717DTOa7YQ4EB[QM]K=DE:RD??DX::@O)_7
AJ+_R?@VAS,L2?CM]NDFHLYIJ2W&&d^BZb=P/OC^^#eEW&]#?UO;)R\#eBAPM;W<
cG8<V0K1>N:4.]cU:GG-3Bc_H).QW,>LK#+P463daHKc<:V??(a4aH).SKBgK16g
._F3Q)+/&-MdQRWF->MMZZb;f.SY4;X>;&BZ[N[QKG2)U+?H1FT#:[OFdO3U-IFc
M;M]dON9&B,0(]8PdX7)f8@V+_TPJN9adg_?a=A05X;VNe4LOP=MHG6#U?=KCF=O
LX.eKcY3/c=d-E^45Ja]>Gg,IB><43e,#0#PBBb(d#CEe:W:9ZI/BDfK]R4SR@Qf
[W0S?94K91;#ZVDDJI)46IK?QdI-<L^ZU,eI[OL09.;N^OP,0_WY4=XBW,4,Gc/W
#LSNI1.4#()QUB2VP\[?H0,XZ(I-\E/E6FC90IT5T-HZW0A5d81VLd[K.f)eZ.b<
61_=RbHRfUeN4&F/&gYS.^F3gR0_Y-NG6PF-WP56/Ba+<6=RGaTeJND<YbBBf\N>
W6D2L:T&eMJFEL-/aD4?;,)T^a)0L3eZ-fLIA:dV.QK2AG,>LYHa4fY?<2M_(HV4
M@B;_PB\8K#/bJR2N@P2A<Ea;1Ec#3\.JAeDHf0TG-@>\A))FP8>PP0N?0#3^&T5
geeO;O];D&&L7[5EY^O.IU.BJM;fb]IeX:)PFW0MRZ1>gPM]PVN0fI(I>](@>Y;Z
ZBJEHP8g&9II.1NEO1-cC\YbgT9Z.M?J<E4-<E008c\^aZ2OZSO^,-X:_O=U]AJO
F>^(8Z,JV?S5GRS2JQQd,9ZLe?1T0b]U7KN)KYPbC-).R^-J0PDHQ(8R@XUV\c+G
7f4?c9+0G75)^Rg8-a-)^:E(>eDF]7B90NAdGDIJN<#dEa.=1JG)dZUYEI(E.:]6
,K9XN:B9fd&9-([DAWI(X.5>Y#EK&A63U?\Pab<dKdHX5a^LO,@WYc@c,FW327F:
.G4EZa0]QH^+C+&O-#37,[.Z0SH;c.]FB_\W=TWcI;9S1@;HUBW[G\OCNOT=]5-2
;T/CbD]A;@(3S>g.5f]DcMKNaDA?I8\Bb?<3(4ScFXH2\+YcVVNObNJ9dEU;8(\A
1Y8VR3c<g?8SK72YDcYIOABB&Z\8df&G+:UHAAag;fS;\^GC.9.A.D2Y9Z.P=5JB
SOT+FCGcK\@c_Y?,#/N1O4NeH,H5CVc,S?77HSX?@e=OEg4[_Y3667Yc\[3(1CK,
fMV9@M=L=+>D.(/7&?V5CD2#,GFAXO=OT@2b,:.DRR(>BGN?E\JF<#f1eN>F>;^\
:PF<O_:H),?IfC>6?BeP&?a+P(b8F1=.Fa/GQ5^_G_0RJ@J&1,Ga.H:UFV-,#QOK
e87J[MJO\NB?(>+83+JTGPNR2Q)_Q94KH8Y#S38-X[C3U9<>LE0ZW[g9KCbOYb#2
5<aI#GWIJ>PP;0K^1_2O-JHA=E?D0ffP6>;dU[N+1(S77^)5(A07>N],32g)F[O7
:cd;eJc\O.0T\I,S#=]C+[A5.S[DJ7#Vf2[?2L/b>=[5-QV\1NO[L0Mg/Q0AY^?P
eV0Q(>eRQ>0NW.Z[JKT/:-ALQVTgGKX0efYHQY86L#W]WQFV_fM>eG_.e,Id<d\+
fV,>1OS2OB=G.ad\8]]6@U+2/(T33>:@dB[S3ICO&\dH^;A0W&HY6S37GT<M@K67
_e3RFUX=a046_G-8D(M(:@7U+>C7E4Y6:4MWg,a6^0@R7G:942W,Q37>AXSK&[d>
[=GTce_K(0FDXRG96[.=.R>N=-Ma@D]]bN;WIM<-:Db6.fMVP0^[aCA[6Fb-e)UR
M8G&1=ACdHD:1S?(f=Vc[F<=Q)FO@VTSbW<81DE)XJ\D3dCXS[B@9YU+CJ@1c&Q,
a3)ZB,,b3bX)G/,=L1CC:A+75YMB9c2<@&F@D;>(24I?(]ZZc^YUL93HI]?f-H[F
LHfKb^4-C.B;[BcDbPFg_2Y^E3M+aXLg/UVUd_RB.BG&_)UV97\1W(_)U=&F9M1_
O#)ZY.<+RU8T_:#:=+MPJ@)c^g&]..PG2IZBeEaeLW(G\8;1ZN-RY;?e2X^/2\C\
Q8FS2-Z?4+T]BHQM7J_OT2:P<641PK\89_+Q7)26Nc?2Pa+9(,[O5[][C+:3gBMP
D.(9>7Df5#Z7HKKTL-B^87?L@L4X36,OZE#TbM][Dc,K<_)UDOQ45:5\&>HWOB+d
1S\b<9F03>,L[UA;cX3.LcS1:[QY8Qe3W6I?C>,Yb//c?<8,X.e1X2G3E<5g.ZBO
FNJ[HFb-QC9UEO2=)1U5^Pa4L#>J6P+R..0Z_3Y5<\)bNZCU+ZIW<DZHT@#a<<5I
d?@]Kd,,_AMYP^(MfZC-[4gCRcJ]</DQ3OSU2JK3VZ]_6[a]>;2(@Y9/[Bc3I/K7
<\;TOO0[;f1W1=fIJ?a=EJKM70FgJNEEN-(D-OfI;@HgV,TA>eJ4T1dE<&R+fUUg
-05,We6K@E4J.0R/&JdYA[0J&R#&\]W698&^\_,Z;V+7:/00?]X.TMBUZ^YTS(9+
)>IU#0GVJGK\YWM&])(d,?/;]&/EcR)0NdAXV?b7+@#.@H;\LcV+QA1c81K1#A):
E3X@E[+,G.e[cV2Xd_7NbYbV#CadW9T,LDJ7Z9T4,a7@UDY;STSI.+V@TE>N\SID
[Pe?H-eSB73FXW6QWfG62^6Z_D0TD,2MM=]T4WW362I1aU@:K&W_WVL:AY[&CNY>
14V,;Y,AY]_?IV72Y_BeaFAP&\(=R/&6L1ID[RJIBUg,H:c6I?BVTR.UVeegMeJ]
.Y]AU6DC<3LT]6X7P6/UX]2]PH;46^F(?I>U1IKFd[/bJP2U6D:.68H>]>&[@WOM
]5I1f++2+;DG<J;b,/LZLd0>H?BbF?,3NSNP]88T_0_[DDB@)FSf8ZPWDVG_gQe@
MG6X^YW2-F[-,4Z;;&\H)eOf7;^UQ2^XP@1J/E]E/)?G9F#ABZ@YRPDSAf&fXY]7
HA4E/DP[0^SRH]&CJ&J(ET<HX+Zb;LK@N,;(DFe>I^XOGP?(]Cfd8@DFHD)-=+4O
QBA4W4JPL6T5X_)2A\_FJKNRA[??_(;^A\V]3?Q_A>/0&4(QLZ>?@U6E2=2H6HcN
M@e83Pb]FCHY/^W@B#;aPGQ;<+J,QIC[eQ^=#W)3CXWXDRLZ_1ZPRVAO/;f-c.OL
[c\A4cOJ7^cA-SZgA&(bSKcZO<6WNSGF5=]?I4XS3eUYZ/2,1;T(Y;(.99Q__P)5
1Y;T\_?S4C]AD[X2E=fe8TU()P(T]&PE@8d>WK_[cf2\_LVI)RK[W=@>5]8W0?^V
Z1U,>,/RMJLS90WeKRM^[?>@C,43c8>f(DF#W@[87OJBOa2:1K,Lf[=<ELd0Y2AS
LB/QR]P:;E)8.[Y2cXHXF+7DM64aI=T;O#FEN[15:#X@JK&8g5(VA-HC6fMVF^V>
(?UFJ@LE?]WeHeaQJQNS[\MdM2:YDZF=H,D=27DBTVgM>P&B5cY(DLU\8gQg5I+Y
VW&<7V(,g6WYS2e/@?^H)UOD\-><<X5?XW2(3^N]Z(KP9S3+f&F8F_<Dc0>J3HM9
RPE2/DJTQ)+/4-Zc]G>FN)9?LIST[d3M+ZAJd5M>JVe0?Jf@,:H;L1eB\>.F,[QU
NKdK(+V(gA,]\O]dR7_QHPV\_]J\()@L<>gRS[XBOQG^#J[5X)_8fS-<e4,,8@M7
BG_683+VO.7(U,Y0R^S]I-+U3Oe/RNfbgc@f2]MX_g:SHbVRXW>WR7eNSA?3e7SL
GAgNYd:dGB6>._KATH=X4X_MFP#WW?#?FJ1]>6SP+CdL=Eb0HIR;a?Od75cH+XDc
Qf(M:6\GLL?^]9/8F8S20X:AfZa;:S2cX4@@D40_3:+3:^ac^<IOIcN^9M7YZDG<
S(g#+Q)T7PQM]CPW9H)QM/@/_(;O2EKc:GRI/\K(LN.CUVc[VG?T]HZf:X@UU\XY
A?;.>QA89#b(5=5?:OEV+ZfG)N_EW3#9SP7_bU)Bb4Qc#IF(D6Q+KB#4_=0DW,H/
+#RC:QX&6[B>&@e#,)@TB6DMC/#N=G,E/,&_E.G2?&XURNS7E@1G#/c4S9;LDC)T
2aIfd@Se_:8CRNGD2gY\+&Z9a)H77S@gFbcUWS^LV_9M,:;8QM)0&Z;2#&fbWU5^
UC^1L<,g3/)ZO[M(e_=<0:5#COcTc\+e8H410Rg_#1HE(O@/BB,B^P5e&0-U:6/=
&H9+AD/1,L8&<,QGQJE(.^120AMEYX58_\6EW^>XL;eHKOSN=_&,XDTCF2/dGEOV
N8?O-_HXV9Y_G3HJ9JW-=I9JWCHR-KIFEf8&#<bS3BIM1=Nf@9,>We6;X\W3ZJE8
daV,UOP^9gLU(JIWGI0K:C-[;&.GH_0BMD=J?ZPf:fU5_KK=RO5?K>_I>\@Q/279
S@HGRYO(HZ))K8XR:c1BfG@0>=6D>JN-9Q[5_#>gC.Uf3b+=@ON5((G:[TYDC0VT
F>7^D;.=&FQ-/-b@7d1U<,[Ae//SbKT\d,cR?YA3AJEI[NY5;+D(Y&J^e>I;EScC
]cDY_X:_7WIYFEG<WLLWBXcUW8f.)aMSSOD=K.b7S2Q&2bbE#6XTYYXBCANCg.+:
0YI[&4&RL3g;Y7]S;BP/DQ8#E7c:,IQgETIIb_^@d:@YJ8>Y<GH/Z67T,1b/SZ3P
c4/0;#Ic5e8<2Z<;+eI0ZeAZg[<2&JIOO?&WX3NP?+&2RULIJ)G0Ea4?a78I^JFV
/)b;3>\=&aGAaLH)SSfgJ73JbP8b\AI,Qb=8YdWOC#@^70<D>.&U(cRK#c&9?_?K
FCd4-7&3&4((QW<R2K4AJO&fH&,6[PRIdR;L8-8Vc69]DZ1RfI6K/G)0/\,G2?@E
WfH6X7HH<YI7B#HL1bF:8RQ.9f0BT)@8TVY?#=RV9PYIE+UR[c<F7VL=/Ha#bg<P
#.L6&4+RT<0W_;2G\[Tf5NA.0OY2eKb:GM8[[2R=;1B^U<5ZMB2B_4#cd)B>4eA[
,gaV-Z0bZFW&5[4HW)-T39-6bL3=H#L]JDR.LQ_^9=/RX&<6X4dI.4aR\,R;@aV6
ZA/B1?ccB8(#3VC-6ZTWX-0V-gg8E=C,97,X<LbMa8O1]PO.4SBg)+QL&T];1a+f
0->_OM=^6ADQ(a.EHZG&9,=-5KJFd+ab-Kf7UB0=(_D297.[[TD=1LEO3:C-+Rbg
AVebSYN#HSNQ/:]9WTOaY)7K\QZS][efS\->YUI]^+&c+O1?Mc+5&]W&WW@2b-H+
eHPL5G#^614aaA98-J=8]\V6VQf].MEf=WD;NIGJNK\P\[0Fb-T:gT2Ka6Z0IT1#
\[/b.JG?A;2</CZ(6)\ZR6I&VIN<bQ>0)CNPJA[WHMa3P-8F^M2E:S_aC[+R2\@E
\47DH#4++]O<TeXP]C(<+;M#?aTK/Z[f4H>+HT>g4QOY[X15fDKF85YM_LWLf<;f
.+D367g@\M,G#X2B+M6G9VbP/3e65<#^:f9-&c<6c&.L)(6a&#6]]NbP24F+JNDJ
#?^A9bLT.ND#KC-5Rg_:+K.K=eZFCM8L2+DSL<BeQ<#(O.2f/@Q0#+&Pf5R?#;DK
:>SDUCMa5&I<fXU47Oe8?R+D3.IR0H5D9.L^5aI;0[TXT?Ec;X-1)dbZP)2ISV62
P58_@E[\I??_3[./M6B^\:?A-3T>9J9Zf)N]f-G[.2VUg/W0JP03)+OH4<8a?R&M
d5>8/d<2-dBPGS[Jb:UN0>9XV6FGBd-NQ3?I1_7IcKRQ+UHM#aP/Bd.)IYHFPe3=
<W[.0JDOg-JJ:^c\BI\aBTTB.FAY=7bcE)8,RH2P.0>&8<>)d+_LX+0<GDJ@Bf25
JZ_(<&gKW\[W9)[DWbCI.C77@K^KG/cOE6.fMa=5(]RN[]b>,YPM5LBUF(eb+U?U
89J8d7\_=L+N1ZR;AZRK;5,Da/Z<.0C-?=#4L375/]DZ?CDZ.VCc[PFV==T-?YXL
5D]9W08BI;=f#RUbg/?gORd31(K8GY<S<FZAZ//?HCBSS#U<XN-2XPgRQEeR^D@<
3B,5Qe/L17T]:a-=LQX[-Gc72#]OAD9g]0OEY./Z(^b8IL:&fF;?0L:/Z>81??cB
-c-MA?9dG::Z1=4TH+W\4\ERDCC89-SMF?HX#KUDU\/)][J,T,eXOQQZF/g=I2/R
72:+B\I/T4,bEX5MF9P=Y(+[+J.)_cI8ND^5;8/E+/J?aB</cYAc@gC7=df_CO;Y
9HLa>^(M1^Ib.^g)2H0]9G0HL(Z4-2HF)H-\[W(CAG[]+H)^e<?;Qc\B_FFA\2=+
_cXJ9QBd\JQZ6FF9VX6IdLP(bYI4G5(<:IM:=O\4Ac\CXQ1H]6>651?#BB<9&DBD
^:96:4&1Z0L@?&>>5L/(,fM-0:?)[C_Q><KK0\;5EcGf4<7^J+SP1?+:<[Qd@X5F
21IZT/5<&>])2E5bYO<>04RO&X.)TAE5;bWUY2NaY7Z5ad0Ta2RLIf4#c/(7=A<]
#(EAL@6b@Ab<f\K3LC946;.;@d^HKT&bSX(8H^^_=TXWI?U5\.Z5L6@WG:#V7g^1
GJO?[TH.)e@X[Lg/W@UD2S^4Ze+.5@:CXc?A-2LE5FMNc7<b<2Q4LLTMaAFQUU,2
1;dGMXL949e;\4CHL3\2]R13&XJKgKB?DY2NK_G]Rc7_2;J&J85QKXWTCQP#,M];
G?_B3cULO5.0V5?WE@WGN+=GYVMK])F8FUX=.1;QfE_f;@511(1W?I<1-O,5Cc,G
M2F/SW3C4NS)N]DQ[XPZ;7H9TP=/L?RGWB=#H2[SVDC0Xa&P6EY5Se;Na?a_WUU@
XLZU8=,a_P9&-66[4CYQNI8WMPE+BMX\7OR1e//>>/M_3WOZBO=P6c]cHGeE&OI9
D>L23D?ON-UF@-GCQ?WOaHVA?MfAKd-W#EF673OD[5c+3;1V0?#OQZ?8e[X&KDG1
W5.Qed,eE^P#:Sc_<OJcAf\[ZY/7g>gFb8J9.DIgQYHX\3a7;dJ3OUZXDef-<gYf
:DB.&+K_JW/CUSYC-P-YST71g=@42WR-e0&-\S3f_J9T^dPRgC^^&M<62(]MT\HZ
9e-K/3VYAJ@BZ.M@ITNEQ3M[>TQCLDI<c#S:S/fIdYFHf70Q4-TEeM0;AT-N),QY
?c7MAG^]gY<9J#&0_;=J1@M(YIe>^W(e.?0Sa2Hd,QSP9T/S_@&[P.Gd+b-Ub_2\
7TCS8\d8[UU6-BV4=MZSUHB0TWZBJ4WZc])RUb#a5NWWBCK<//-R,W>>WJU1U9a-
I9;D?C_BbQTC[&NT0gW:aW2^M72+OUT4GO5E=c065OdKd1e;,?Yc6-cEB#;WcV)]
GdV-)6XU3c9TK/V+eObZd_YMa+HN;d=KadF<K.:0LE9:Rf=2\9RB/aRS5IfH)SaO
OEF46)b,g@8JFafcIAHZ<FVd70O72LK2M[gDW1T7@G2_WJY5Z+1d,Ye7U]f&Pd6C
1Y]R8]>bga??f3.f(U(8-GUFD=TW.G68bSd@^g;fL>A<8<#5_f-KATWc.8F9_bGF
>S.,GcL>8<#5;UKY0LG9UY,+1--_(Ab@.2EXONC[9e7b.a\X-dW7R2-V<bR(/MB&
\-BR7;@]Cc/8I)NF7]aAWRg]bY?4gW1U0MJ<Q&)PS+4=gAbL&BdRg.IBL<COC&11
)NI/DB-B-63T\LBVH,5;HJ<>)V,J;L><7TQNgAG,X.g4&f.GS0)UO&NdC;700;^5
KO:;-K)M5>ba#>f<7Y@#aAE_SX&ca\E,WLA96af(=#XP<CG/c6&bK,G[\][_M0<g
634@aD.4FfdUc#N&P,W<EY=2J,@E_(IATdIXE=J?@R6A+)W(R?W/EL7^,,-(\@(]
#=gI^2NLbRB=0)e7bb,<0@K8F_&ER9^QM4M?^AB2?WYcF>QaI[7<CCISS_bLK=I2
89-VC?[NY\gW:<#[01gD((TS^-PE[JeGKZYNPS#42+<M1I,4?DB:G[@SE>[,H>Se
W>3_]:9+0U9:@TRS61OYH&+IS6K+)B;ZRc(^TR\,Q6;C.gS+__4aZdJ>[(#29Q7N
CN51G#C-10TKCA\H9TMTSc:D#@M9dYD)@dc\;GfE7<@@Y>M[C24e^4f^XY:UdF4)
<54_6ccA;-/]M)9&]V44\C36MI;9eZ#B5YMTdEPT00bI3UFa)b9@63/9E475Ve=f
2d>1YaPf:7FKMfK/,Z2V6=EY-TI#DcFC[Z;\e.fYGc=dWG6.Y>>:AWL39A=:1+^N
L<>+?)6,IG[Eb<R/S[]BP#@3b=1O>U9#E<]TU5V.]-Z>L9O<6TaE]8a829D.#^I;
fM6+=M]B:=RS:4#RV3569VRK]UU>Y;U<);WaR88[?&WaZ\97FXES;>4P&fGS[P+c
VY]A8Y3]1/6c#Bg,6^F[N-[R3[]X#0]GXCW+f\9.3eZJLLHUHAc9>b1@9.TLLY6f
SZ\)BWQ.MM^e6Zd7fMN)GJ:B>G&YOX.55O&),:]\7DSX)LUIN7WQePXV0N9J4(^G
@&PbB)SKMdWGXLKLaa7>(ag7(B-1J(C_RUO0ZINg31,+bX^=3:5\aX?I=Z6D.,<G
b[Sa<TQ4N+)Z=dCMJd:fYSMPL3bR:fS&K)ed#;3^gZR=_U>-DUNbLCXdRY43B<EB
JBVP)L+,T97Q013F[G13O#e9KYL;QL&JFO0V&X\M;Kf?7Q3WY4GB+<O&4Db[KTL>
d5@XB+;<[?0@0]0Q3J7#[>,3g<@K+?fB6LW^<Z9;,a6KR.S/Tb_.C2Q@?8G^HD<<
_X_Z_088d-4T]MG[_9fV4(]2[(g8QH]1c=;?d84ce4&DKVA45@7c<5H\])T-Qc1O
X8.@(-?A^Y\62a<;c3(QI9YV3FdDg)1Qb#@Y]?\JDb=]@UWG@5K?N?0-4#bC>->_
\/Fd6D5T(JQC\cI#356#)M<eP25fTK6QeV3S,5.76WHEHR?B8Z)@C@R&HSM(6ITN
cdBN?W@9:_MPgDXME84PQ,C1:eK,YLXAMV>:I7cP_7[II(,#P^5(TOS#;[3G>bX,
3EG4cHD?EVYYe1c]e^-JF+;3_(<cDMYVc774ge0@eN>RIO\64)[450M>[641d:1=
T8^;7\VNbK\F(3cOVZU\5(,#,-4dYRT2\MbaQ9F=P^c&g)f<eP&=SeT/2R:SN71;
THg76KGR\9C.OM,9)&,4dfH[2<90Xe8I2(gMX](TOdH;gTK=[e6@HHL,[0.XM/)c
NY9IRb8-\(D1;0d;S4(Z]]:K\LO=7:0S\/_dQINKB;)8^3:f7=e38&PE=12?gdYD
YJg7S&-gVZV1<-9J_#4f.=RKQ7[QfARS_7:4Z\fZ1QKgf4Sf;-&<gD2UZ^JTJXZ7
/cQ)eLNOe<d^N=O2N_-fRf&Xe2O)RX=7PDc\ab/(K)4ge(6e1FfMX^^[\?Z9eS\]
WSXCQDX;RO-X4#(P+a,K#^0ERU7Lc8^^P99TGFV0aeHVO,46C)8IW>P1AM]D9>]]
ZBa)TV9@g-C=-EB^S0M(F7R-[/[5fM<AM8VU#\HQUG^bcE6R&)@3R&VTBNL_L-./
007)N\66I,Eb54L51gXFD?eUH5V^#fR9&]Z0M8#_QYGPGgQeO_Pa4.1eeH4gAO6_
c?WF^=fY+;?W]5>?D@H=f@])A9Eg2W+QIafO+FK)T23@/^S>:^IY.2IX7RCbd(A\
0G\Gf206@H<e,?aRRKa\+@c6Z=1F01a;.d^7]@)S2<PNV4)daS=6^UK]+L)IT_La
8N_#7Ja(\[Q?PF-@)D7GB4W^-4[&LdX6fHHFL[#daQLC[ag>[KY=/6J>[NLa=Oa]
_;>B<gSW+:fVC[-&2Q?0)M:UR@Z21S^;<O9OG[b5@GR7gdff(OW-S=1D9B_Xb.>F
AJ0,<8YT?:a4IAGZ@Z:<Z7ddTQKRJ8:c@cg5(EFB;I:,<]7;9J0X1dU=56,DK5I(
[VPIJDYOAS33f-<.7FB#YAIEE;V9)\O7:a9VHffX/&:/NMCYgQDQLd:ZCBGC2\]Z
H#RK.S\Me1e<V0LWa0@<d6I^Ne,5QaRD<I3HB:Z8-eCW-_;<)7(c^:-(RdE.C>)V
9NV,=<8P=9&3GOTZ]MGMAQ;2I,OT)<V=/P]4Q5HB](&V=,=A1QV74@eN3[FBIOg[
bN19eADO)=P?4F>^)^28QSSMg:TdAVKG,PQG#a#<T=9@W817/a5;#UGc@QFHO;RJ
#&9_O):F5XA?,&G=PJ>18fcCG::,.&FgJ6\aDOB)bU,)4aI8g)a0e1S\.C>e;T2d
QIe\bQM#]WcBB6KLM>8RWbFGN9EeV@[EKZ9)1AW+a.9b]?eaZHLDN8Jc,74_a350
2K6dD>X#SRMGb3#]+#49UG;[C(2T0V/Bg)EeBc[)9/N.#3cI6eYaceKUdLLR3_d@
&Me:a4g1T_aP9\^)g_#F#Gd0]PE=)+d&SEe6\92PX(I@d\5^IaWJ.=[_D4O5#bSV
CP;g^,K5V+>GIOXcJ@e:e4DU:0@43:714B_WO_0#\/eGV9)_:+Dg<CYR>_,XMWB8
.=H72DMMHe]T(9?V2ON0T1[\e_FeUBY&fd[bAS_a)^,8M3.8GB3T->g/MZ/ZRaQP
PZJQ&?G8HOOGSPW?N7<,#1QJWX5>Jf-FZSH_T5Agc(HK=g;GBS.<6_^0M<2TFSD[
XCbR)1H99dL.#94_^&YA[HOe1-f-YVF#[&B6Lf4LdZcgDb[\-E,6[XHX8RFeMacK
W3[3PK_7677NMI886T>7=(S)](X(9H-.@HW2,Z7#:)g1=Mf>_?1B.b/M>aTCPcZH
f=A;;E_+A)PP(7<&Q+H?:g.#TP@?:QT5H9Z;a=4g#1N7-P/PF_T_Bf+_]aVTS>&7
#;4a#3C99OUgS24G?\&gDcYJL4=Z<@a-WIIb(QPJQ78BFA8_27/<Q<]4)eJ8Q_<W
T\VZ=C>&U#B3:OEWWCCE0V.LVE9J\U--U+X=.U8T,-WCdTH)4\B5A\COfF+S7?Ug
4#EUW5:ORFZ2HBgV5?@DS1W#QfRK&IcK@E@:)M4G5<L&811YH[-gD?/#@R-)GF]A
1D81GDQQUYW)526-?+Q;G3b5J+3=9#=a74P+RG]R(X:<:>:>,8.6)A)]B_LBU4;0
bXdC3EZO39^?B#[E)BD26\Z92]L/0F#(eTBNS,EKEb\4;CfQ)X[cB&3CP@Q)TPGK
)9:<FFD258d4C.=Kg/..^S8cBG[H3e\S,&a58(0=WJ&?af-15;S\2[V0#LV9Y81R
-,G3+5W9K7ba7?+-H5Ua9PN27V)W5cbAE<GQ7VG,H91,_)0T/aHIc3d@MHSPeAFS
&7KY[:J42K@CIV:Y4?9V\TXVSU:UBTP5>Na:[b>-]B@,&_M7&MG:R4LY_HCE?465
2g)>#LKLT5IDF_L;O9AY<SR<IN]1PdOLZ1FUfd(DY;8/GfTD]P0T7FV1SR^/Z[>b
QD]L#0E>I=S2M1O:DNG)_YHL#[W2Yac?+GZ,BKFG4aU_TA9KPcf-F@9QO3da1-[8
VK(GUH(P;<c&ee:4M0=Eg,fc>&G/cbBJE0e7YR&KH]\(S<L&ZMHCLBe=AC(EP/3R
IgAc\8:N:(<2e)KQcLPF(eH[g287CWG88L\<?)cAb+UN.V&2S@\dg>L\>49F1@J1
W,[^4:&B6ef&dV80_Y1\Q@ZgTZIJ8@^\>PR3GdZ\Nfe>7[[CR=f[ON[V89FI,I/C
UU[<7HNTXQ)=]&[^ZNS5G_>?J]4IV1)GG;J-UTdX<@=M9#;Y>MK@2g00XEZIg#/P
[R;N^;@\g7@=_0\7]6YR^JL&QA#^LG_XU(KVHH+7PL=/CPHEe:(_@fYF;W[@g-Z=
TZ@QMTC<>61JI@#42.I3]K^,Y3Ed+0-J=\g7W>P+ZA>U,gR>eJ=JL7.aG-dEeN09
R,,Xf[LED+X43&/[ZK-Z4X.BbE>8)8)fQHU//B3L.J-BW5?8)\P?gg?gB\L)7;V]
4OfCTFI2O^4f-1WX#eV(R_6#RH5^-XJ\1d(+<_/L@]U6b4;g?aK&]DHL^gD2O)N2
dOd^<[.<,O,6/]DLFIQ0A0>S5N^[#N3d1=:gZ6g7?T,UQ8KEWJ&SJ(YO/:_MK;OS
MMOD7SA<+A>K8DY^[_WF]gM4.]>1E,]@)]UF)F58TbDQLH:F8,Y3.38fb[?02RcG
]R+TF[H)0X#XXHeJ,EFceU[I>(MH-#F@8N&7D)K60,d>#B8A-#TSTA<&CY<S2AcW
dXV\P^/TASKU^+>]I08cZ8KRFA2GM2=-c-B5NEMf.4c<\,8ZZ9O#Z9\M>,fAFefe
OMSTcN.TR\aQ=>a?7<EdI^,]?SJV9c^TeJ3a63&MgIDIKZMK+0D+[7;I0<TL:-XJ
=aK#76=GJ/CLWXG:(SB&N3[2Q^8(,#NVaKHS5=[7,KZ9,c4W4C@+9MK)B0K+)89:
VB.VO1Z?Z9Xa(RU7RdT/Qb1Y\=a?<I:#[BG4O)>M\bb?Aa]LMX3SX6@MLZK,PBR;
0WKU)9\^=;+KRBVYY9RLZV:L-)M\VBTW<[K=W;Z\aG>Bf@eJK?22]cQ5We(8YXVR
bXB426/_K2b=fSMAGSH99eD55((O\,M0_8b_e\aQ&-\X;2b[fU4?W>b[bGfPd02&
2+S05Y4ACOJ()^:O@>8IG/=S@DJZYU+Z;.5DMZ90A\NF<gDH2]K/=4[&-_d9X5^6
Ie3P&bZLFS3/(X>H0bCZ)[(+PA8,(dEb6F/Q18\L-_QN_@O)ND_VA=QLa36/6NF]
0M+C)J/HL/Q]MJC/-)/O\B9G^Ea.O)fFBf299C9eU6[R0/JVP?6&6HF:]N519a?^
Jd7<3b2.SJ9Ve]EGNK#,E89,VAE_7>Bda4);DJJ4\G9HA/RXZM9HY(454,#5aX\-
^C#X9Q8KI8DW4Jd#FFCd\M)7365;JT.JU;T<=3^f+DcI>CeND0DS;G2V@]]QfK/^
XMSJ5Y@W6H(#B/58fZIG;1ea/PG#@FZD3-JB.C=ZHEP3Z(\ZVRKf8+FeOY<6W4&f
N+8OBZP<[8TdQACO+QT910YPg&->&1.20#79Y)R3]R-e)e1#37YS(Zfa_:U^b4+N
,+)C5@PeFCf?I2E41H0/(NN/;I7YH\G#1+P#I@8Y3UVY/+dSWf:^88JZ[37?2@ZI
7c]I\:\eE-Y1:R#),\[#VeeC0;6bIAFJBb9P=B[+/@]UHO6c77[R8C@GX4S_<H@,
7[9abU0&T[3^>ScMCL6>fLO=G:6aCZdgWCG>Z,Q8TPWc+=0+bGUSMT]e46]V.5OZ
5)_42\XZ/a/-Q,=P,BE]K^[g.[-faD^U>19fA1eJMN>BJbMbP/8OR40WS]_-ec<?
_>#ETEcWZA9,@P^0DQ6=4&#>L4V,TdD0^@7I_-K\NBHa@c3,9#->2HQ-bXUKI,F&
,?g_KXI/bT6/COFG8P=OWQ])MUaeM,^NOLZC=?>KPP.AMg8\]:cFOV):1W6,Tge/
.=6+/FTLZBef8?[0.YZ<)e8R\>X5B,H,KUD;a\_2LP#]a>R^3H#;D@3OWY4[WZEW
>[N.&fPP:T#^NK58f2^YIXO.G^7#73?43J<O.3-^]-ZS_XPY/G\]R12eU&MP7N57
X2)W#,_5\OfRHZ(CC,b@#-O(D.]+de5=]O^_aDA>O9R[TH:-cE9(;&Q\ZY#2YKC<
cQ:V6N.IX4N.2c,c46EKacAZeBE3K1a.&B=[QP+7/Y/IE:O8UCRA@(2;gLTGGRFL
4\S8NO04>^C:7?JMe-VTd<HE>JV43cVN@E9g1CGd^)T-.J.VZfH:cTXc/-gY3>#1
,-\8K3IML#GOX:W<\M9#QW-Sg+CND;_H2bK.?&65QLfJA)9bd,\JgE<=f,7bDX_D
YB3ReAU2U6AU)#c5HcBMCLNK0:\XER4:GEQ@KXN3a/b7(L15@8efIGW)#<JMSaH>
dDZ8=+T?FY/,FLQ<W#/V;XW)^(dVVXaBD3M]E/^Q(1L:g1<(CB^Z6Pb-]9eb_^Ee
?eF@T83b?G]<-NJ3P62K/S)Y;W6.;:EBS=3P]cMf]bBab?XYY\YP[[SGeZ#5-Q>G
PG:R,T6>M;W6UMc=+-GbV=X^#&^6A;TH=M[RIcCEWQ;#([S#c<6#Ye(K&e#T+FZ@
?83F;X?8>J[\/SAVE[B<TW&;IU5d9O;#gEENO\^SC:LMW^T2/&g768SCc:BcA.//
4Q3:_EgW+W9dI4EPN;d)&[FEg#c&g(0E(,>23K/)Ddg9b0]0_=g_EdKI#,:Y/WT)
2\A9b?>MY[Y_CRf0T]0edG-e(3.+W&F>N,H=N2&NGQFeOM=A,SV;AFC8B/:TJH4N
O\9+K0[>X3^.UI1OS#bOL<57RT:Nd>V=d&\a&]_XT90/.32M>6,;+FdJ3]T]5AU.
XYXRgdGf[b.RS=+Yc7Kc1SP\RP\:D3C;_ISTOP?\6_^[A@JXR>FN&.QDNP1Y&I;-
+&2:]Y_#EE#@(A]IICK6_,Q?9L>DM;PV1-M#CfY0KC#4M1(H>+&,OUfg([d#W<:g
^ZP2)7Wd@UE=UBJB/OeccO[(X;eAH<=F\8aUDZS7AJ:,5XZ2g\.>1Y:S90X+X;=0
+<1dfKTZ\,7<JMAQTJ0:N\9V&0<ALG&D_3/2]#Sb/5L?.a)B_F\f8MBI5d.3,9,<
\SLFXKe0H\@;A#P@R[S@b]1aJd-8C5Y/)4?P^_=N(\E5fVA4-V@,PB\:3EMU_aQ[
.gd#7C>@4?8ZNZVF1-+8fK.X;Vf(ZWA6(2T([^/7GeGGGXDgbL;5,(SQU\..:a&L
@S2a1aVRF^ccI=A#A3fG2EP+FdK>)]R8=7c2#VVU@IW<BDa&G=C9.8R=N,M+TMEU
B42VV95/&1(dX?a.7K;B\/:#a([(@&_EZ9(2G<4DdKK[<A6=+B@P,XI;(L7:@gX9
g1;_>D[UMF&.Y@IX5&MU=/LMZe+AE,2Z,X<8-)IK9cKB<Y[:Q<[a_Ze)7MdWfI6?
[AGb.cdZ<V:=a3Jd=TL.K4R-EGS,e96DBV:#RMUZ?RfE#:O873,41@7c<HMX+D[e
5fbbGJ\?50SRHTHX9-Jc+P61gU\bdP8))_e-124gK@_7.>d&Y4B.cZS=?&&K([TF
gZ@N+d?(5cU^3>1S:.]_A?6^MR&1d[;XY)VT>RZ]DS?\g7S,,#OA?V=94NTLYSR(
b7Ke1.1TGF?73R=NVVG=G^WA<c+(/3S4,A=<)O3Z]c184T&1W?V84;JS?M/?[UWd
^Z<&LS(;]d&&_-C-fZa9&[/HR&CU&P[aBGJY5B@]Za=Ug[T@d[J6cY9f<g]]d,_3
=gY[N#1eASF.9&6)JT9>Z#bN8BgC;>]gbOFL8P^-O,#Y.@=AN<#S\M3Kc3=e@;G>
;WKdX>J,LS]6A0[M5Vc71ee]J<CWZ3(.c6+^Z>5FBfL0QT]]Q\176RM[G6EIObCb
eKZZ,7ZL/\bC.\T2Q>PW#KA_C6WdQK>U_,:FTI\VV@c?_UZ846=NDSeI#b/dI,,g
6MKSA:7-V[Yg2c;TE)Y2^2bF155-^Q(4TMcZa390:TXd6FBBSB,OcHM6R>8+REK&
4JOQa5IWU2B5/X=_9T&]0>FUHbe&2)e?BFR/5]QM9\?6_c6(E(O]K&57)1cO(@)Z
.cQD:,>)Ud(CQ:e9Q/gFIa29]:X]B&3d:.JK2e920LY&b=8HZQS(C0EEd^-R)_0:
.BEb+L)A6(FbZU)7d\@EHH9KU^P:#32A,/[8/K<SB&1,/0\gH5N3I_cM[F(;7#-P
Q19d95>G-H>e9+>U)UfcCg)VB+1W_K<QT,IJ@M9,CNJ/(=XZ3dHYRFfW\.gM_Rd1
WHIJ29V8I0fR\]\3/OEJ(NATFc,D-VH4^2=W^/)WX01&4<E;1^?5E&50[X:&_XD<
Kg17L76ZDa7LF8N3fTb=2f025YYH;a2LcT;c&KG/Ua\YF832AKU/0\^6,GX:</5a
HAb[]OHG>KK2,1GT)G@>;>2S@MGOZ_TfaS.P,N3BMeEM+I1#N7R<0C6Q4IJP5ba=
+QF[+IJJK<aee(FF>7REOaU<,&?4I02(Z4:A&(8G7gW067c?3gY[#.Z6KcP4ZDN9
1)^?]1K_LX7V2(]K/#5FgbE]g/X5Q+6g2WDLUS0(#L4dN.XJA&R[aN]T?BK>1DM@
G,>+b]M,c_QN37Q2]X1H[@\-7.?e-bM#@M^[X<;Z#&<A9U;>5^f)+2Q.LQP&KY]8
BbNd&J:]Se1O-G9EcC(CNQC]-7?6.Ta1e^C\Z@U/[O#WKQR@RO]W^\FH9Z.=]>OK
W5+7EJ3>[cO[&./eWAUC3,5&[b:;9ZgF5&8cF5_9Z(b9&\eH7^P?(TB3P)a1VHXW
L(=JDW8eg=DIX6f7WGb4:J9;\.8;3e4:^LDXSV2(Sd.c/PX[9A?=S7DJ7=TZN75X
);^T78B=L:GT?.TfDL:^B<aQ1?2-B^:/=>ITB&a:ETL:fKD#@+2&?\CO:d&.A0f9
8UX:_<>QK)_(3MH5T^)JU&9).c\f#=)C+7G1SUF9e7]-OB>5&Me(+-F-7_BW],Q>
M.&R(bI#VPQ@R.=7+JGg;&LIDT:3:8RcbZ<ECc)ZPS4J1>EVeQ\F#8da()=SGJKW
,X[98?1A0MdN8+Xe/\f@\89&L-O.R7+6.1#D5YIZ^P>W5ED06M@Wa:JM<U1:-D@(
fE9.M6306DR,;2>GB5R)30>&/7D?P9@&[f9^XZ[T6BG&eGag>.ZI;AG1dF0ML(Aa
6:D)9<<a&LQN+(EIaCfR=H,,S#DH#)>a@8aK-N);,BXZ+:fXI4J(&\_TV7b5&#PJ
566WXAGTg^_d1K_CSKe=7dB\A#F(=5?8];=9;6Sda45\J=NY3\FDC30X=B_]&ESA
>MIB?bcQ,:BVE(B=#;;VRL]K[f/+SMHA<2c9+X4-:^7.<5XV>[]X,A6\;/\IH(]Y
YV3MQ)ec#a\Kb.,0A+0_@I.GQ;07e=8NOV:)2:A,b>OSS+E-0.:=-MgP9QISW1YX
#SG:L_B;b:S=:XBT8J1/8#AYM+//H6c[0[EX+Ra:f@K9Y8E(KSJf3b.F9GFBcWWO
HBH23/c]8>LB#/809T)F#YZG,Y7fG@Fa)3Ic@\F66NAF5,ad)eZWOZ>TJ)dEP<.9
V0#a&IQP)Y\U,KO^:c6M9EJe&K&e./F&eaa=Aa1e4PF_GS)K=?.3<;R?(2<@_=W?
FU5^BT_5MRC^b<b53AFA:B=+.:G.)V),5Bf93Kc]DNRG(,^[Sf/G\O9K1H3Y39[1
4/MSIY+gUQY:UbGIFUL0TGN8#;D([<;U:DB=0VL3KF\UC-C32eM>.1^PEY:BPT+=
787@I9<a;P^[#-W62f5:><M5)DI\4P8UDaQX(<_[PU?&+5FU&KRKLOT7#Z&@<0eF
f2MG_KaY<Q2P1FJI/MaMUS<)\]dT<-bLMD/D?AB3N6[MSZ/]EQRRO72UFD]J.ge0
/G4&>e/;B\TSJ9A]=I&9ZC16^:<+/-=a2c;>>+IB@(6G>A+>(d;7,<838VaLEMYf
H&X,X9DZ6XNW]ZKC:_NN-D\YUQ-C^.(ER\@05(U7]2BFS;;.SQ]&M4YBDSWK^G@S
#P9\HD,T5W2ZbO=N</b^H1-:=:ce:W4?HIPHI1C0\(\ONOCacMVL>N4cgQ_0H.V_
bUcQ3V#RBGC7&>I[(bE,R_<V7N)F58R@/EQRCPPE2R,GZ]V.J4T^F(;X@&ZH1ATA
>^&L^?=G+c\/+Q++A<0R(+U6SCO(g6f^]6SO,)VPOH&@@(A<<E:UCHXQ1^EGT(<Q
IYZ5HN(C1;BN:cNcHeEb&Z=81PS)=CCNHW,<NT[\JA\gKa#T#@?C7Y#4I\YT,TH?
M)QfR[HNRgeC5R_0KH]Q#DW97-4VT(5=;HKcR_c2FgSDD<[4IK[FRP,FT>CK0U;K
+<563O.#M]?9Me,UGZ#e>1+(D(W,9D0F,SZ.3<=fc>BJd:Z:Q:,d@6@W-AH5QgOQ
>3\X,F89;<\L[UcF[M\;61[SXaSC95P2O=\-f1RZWQ.@C-ZfB&/-bD98g]267<HB
2FWC_ETKgX&K/G/P1<#X(,F6a#Q8,0;?gZfR[6UQ#Ze9@b;cX>Y<Q7?9f-1RH?AQ
MS+]UE#f&]M.&\K/O-TN,TaG51YdZ>(.?(T6aZ0(]\DRb]9]d.?+0_dWD_7A^.&Q
bRPgXY_gKJ])-O<&5+Q0G/JX.EE2H=48V<8T0^&+J^8#BgdC[d.VRUWf#7PWfGLg
:@9QUg:I&,NXZ5;MD-]AaYfU&A@>6>1]e@AP@\HXT6b4JB5b@bIP<2eAY<c,>BLc
E\cMS,5Mg[aE]7RP]2ESADW:Q,XXNaaCT\a1Y^M<V4K0M.C_](]4,:,,g()\V,[f
_:]cgK6]^W=WVS;772g+=YH_4T=86YBRK4-_-1_ES11,c)&-[J?,I3ca3ZFC(FNQ
PPC7?.+\?Cd.eSY0Y;JRKf@(<+^)f,9(6NZfJJ[,?VPIA]^HQefc+4(\JfY(5OWZ
4JJNTa[/1Y)Z0_<\d8A70OGG3<-,TE_2T(6/\c,C<EGOb:_HB6>+gF?>ZNMcIXR)
4O9)(#R]#+=GSbWb^D/d2/<cT713I4N5WGVP09YU2I7153f85R7UfP&FHZWJD<:g
-LEbJ?-CO<&VdMYF9U_cJR)R)&c5MF<a/(OSC-XBBV@O-,,@,<+6Cfe/f\aL@N\7
d/SG(Q8.:<3^#\TH,4GLPQW[6We.AR30LZe+L:3PP=#W>V8#=O;[V?baDP8>^.HD
e&Ig1BJ09L#AEVK8_D>^GN4cZ+RTd?()8\I-M#&JPe3Ba[QR6d_]JAYa<,C,5HLP
N<E4:8cXVA_VDK0Z_Be#fYZNT2B7>\R:37KJD=7c_)Lb[?)J9E=J4aUSIA41&DeP
b<[#DG1\NYZPA@8^1J2S2\15BggM_5)R-<-3?^b.\<3;a2ED=LSND2@4aSRW:ISR
Ye+8C#KaC;WJg4UO;P30VdK70>D,&bffITQUI_DDER./^H)_=Be<[:b2Ta8]d]TL
\H6.,B8d./fa&g6>J@5<YGd&5cNa(=K&e>:)EeX767(XJ7=&ce@XaY4KaDV2fES9
I[>\<3Y6VS<P02>6<+YE?2;.W.2P3X4g&?Q:I/?5V2OCP6a)Q1:]V9/:DU=b(#Y?
G)66T>aQL?,dK53gF=4Y&Ka3U6J&f7L4\HF>;VaJNZJP+<)T>-YR)+VBWgF@SJEH
dAIHK1>HR_F:a:H[CTGR[agXa.c15WM@KDfV>LVHHI^D;#@[c+&f9JSVJ4Dd0FAg
9c.J-dfJ?/0RH>KcYX@X\X2P_F]S[/aG&M-OM,E>OE&>JN.,9;C:.N)ceVcU1V/S
)LBU/>+NYE5f<f[]C_e7(S;+e3ReDJCA-eUF&D0FJ(\1I2Tc6(6aXPe,g6)5R5eK
ZGBW1bP-?7@1N.caN[Y.T3HRH-?U7U.OQ#73Q5K=Qb/4P\A)@;4KP+[a1Wg8,^b0
@I6b)./c7RAYS6-16geD[\17>=f0V:M?b-@f,,CWaeC+VH;R>SPa^P9<e3B_B@Q>
2],#5E4.)HZa2.I_)eX.f_\;M?GD41W@f)8XNW>dW;076)W6,VO7XEJ6KSH06EV;
Obb7(2JV4N4B&ZK3FR6W2B66A/?-93&I[;K.RTO7YA1T0J,,Y>5)[0ZN(CgaGgb;
D4/OX/SN^?()(fd/DU>:<ZL9,S.>(0?cW=:QdIEF,UU#YAQc9JI3?g4_,B+f4?:5
8@T0J8^PV6\4(BVW/9)1>a1+#-^3R>19/:f5WA(#fG:QTKa&+#S7+M((@XQ]O=6Y
7R]dQAVP&P@7[OGO-806.&E3e/(<5HN.?L@AJ_HVL8KVRHB^KJ@))S,/+NHSMMV?
3^J]UGe.b,OEU-V@K7890?<O]FcVObWJ_LV,P(b5gZ99E&V,cJ\,_V^)-8975f#9
ATK83.W\@Z#S\OU\W5E^6U+9@\>SgN/N;W92^9-P1.8L@#R_U@#EeR=7#F?g=UZ+
CNf9Ka;B#b561MA@7MN0X(&7X-g--JC<\8/5K?H6<[P)\2;PT-[XdcK\RQ/>OX.)
?OS[8I2.eJF,<ZKBIGZdOG.PR#bddd/<2)9A9(@D-d)@V3ON-.A@WT9)OB1YV0:^
LG>g@J293f[E(EJHFD7HM7IDW:G8<WT4:NW9J>E7)ACbDGP?29c9)++45.B5.@YM
S3-5(&75)dIR20<cB&eX_Y(T75UJa_[DSeUE_=&LXUYDC=aSQGY?5&a:/<YbE0LA
54U:@40VVZeLB,\MdXTC0/B1H?7KS(ZC>(HMOG(?2,e5RJ@[;ZA/2-b\9(VU^ALS
\PcWSB\U?AU5DX.Oaba#0M6#?\DBJZGecM9936?WN35(-BHLRY7,0N6)E]3.(#Wc
04X]PGZadO/S(>&B5b/9O[[/aLQ;We?EL,R:ISaHOcH8P7T]0>4A;OUbK](XAQ,c
M:N@X#T&c0fG6e?f_;b;aAIIc6+\8g0PM^_8[<\NdD28-XEY5?)ffY-B1P#4<c><
>b-cY#JgGfYVHf@gSB,/HGS=>c\Ee:FD\T)-JfRHA]^A5LXIL5^_JGcGgWV05_H^
3NJ^/GEFfc.+Cc;3#97UWIaeM0Ffd[L7bCOd@1KNRa#CEbW]=/C_Pa[ET7fTA&GX
MQDB<H^2]G1I7_U^fH[4H3V:GH:++)_aGda?EI>?>DD]W.R>/L#&RJ/bS]>0U;;-
=IK:P#M.QS0<25APfEddWYA:G,T,3C8afOJD5fTP:PbIE#E.eMc17ZT70Q20P&K;
M&Ne[MK5A/]\O_QOa,RJ,R3[YGZa5QOH\B+7TR5aW9c2+Aa(c1F&>:?KM,>&=^@I
>=-+?<+PAF.:?JB]MH?PEZE4>f5OD2-;YO@YCP_U.-697\<V^Q.0eR8E\[e0c5O6
-G)R@a30X_WM(_FL0U?OX[3VNG:&5a&9)N<4JN?J2C^BOfOU6>e,a>_,^#[fJPP@
>SCJ4R]g29QZ)SJ0(9@R2A#@B;L5Z?3DO3C1Nb#eAI#AcFcX)9=>XM[\SAKK^I8#
F;N=F6<#CC1&4IK4a,0.gV\dU8>G=8(0YV-&TQPAC\6,T<;bCcQcA\MFD+I/RW>a
63WHPQ]KVeaOW727NCTJ@:34g=T4F1<_4Q:,C2SMW9:24K[FZ,+V87)+COKZCBe&
McWV;J:e3F]H5GJ5c=4?(g<\bZFD-M(3bg(,).YM/.)]@?GLV;2)I7XQGAdg7&[<
P]A>FS6TSa(<GP(J7-E@Yf17/J2&W[E(KfZ0Q-9;>>Y=<YfWId+6@7:W>3I6OH84
G4C-_NQWed2G^/#6ZcE:2D.LgGegc(4baeESRR+1?D8N650Q4-e&dGSf,_8,1B7G
A^\IYSTP><2)gWR-dM:&K8CI+955O@P[(_\f>O)NQBMgM>YIaef88AZVE)=_0=;3
_UI99901^IQL>N,O;8FB]5MC@3GGROND[:#(I@,aaXOWXYd\1T<S[.d]P/Y?/IM_
]/P&78+IJ&9Z^^-:]+GI55JX+#]]>>@1\&>]506F9IF-HZSX8;ERO-d:7PK-9]UY
,,e\3b^XS:?TI6HW:^TO?QbY#8;Yf6:aZ#S17.e7B@,/1efTQ1:=5ZaX_/\:U-e4
(I>0VK(e.c3]D(LZfNP#Sgbb<CBV>S@eUJ1V6X+4PBa(\.#Lf7OE?(e7_]5<>f-f
I#B)-d[2PWJcA-8dR=F-P5TE?-W/cU)8ZRfa+K;@SX.?/&4;MC00[\cX<bPP.G_.
gI[7K2B373L2NR)=BIeALI,@)>(S7Z-UC\96-dC=\(/eabRUXE0>LgVb38+Sb>@J
00]8P,cA>5AF/P<8L?HT[OVY.f3&R[M:SBVD2)#R).eb\fg9=JT-+Ff]eI)UWbLF
.O>fR21J2OUO1DeC?gBg0RMd=2E[-\d]BFaBM2T4J+=Lf:0T)G2\fP(RWI(/?8PD
#,)1:Oc7AJF&63=:#7P<L#,K^5KYbc<UW:#1XJaGFY<L^MVF\<IBS?MG40:6PE]#
O3S#&7F^K4F1<86TUOU)<:bX68:3c/X8Wf2<1679Q)C#FBR3A>cZ=X8PUH2&&gW6
N-_HWRTAgR:#&IF0U=8,-MD]:fF\A@L/#:_U09Tg;dD&9^0c^;L28?PfCa<)J)/+
Y:P02Oga7TE^eNN5@/=?Pca)(RdJ)VSCG:XUQ/SA0B&L_c-0.?[5-K/>(GE&2FbB
KdQLO&E,+b=QA_\)?HaT@:.42;@^G8SZ9\(+94@D4:6S#UJ2J9e(8H80[UF_&4<@
:ceBf(7(\/3c4cF+;&:>]aOf0.8:)F#YMI&RG:)FfVF<eR7/b[\&gW/THF=0IM-;
bd^B1X83BFX]Bc=[H)TO?JOYeWN)^O5PgU@((?Ag#4c^[;KD>4T>Td_2@O/C<H<_
EE<<:B1g@S^;ED2>VH6(Z871bLZ<X/F/EUe_f#\D;@[(S^dWCX615YA^9@0PaJJ_
9bEY?Y&B&]J0=M&U>MAFIVN4f&,5ZNSPBTdeFfJ9T;]3g^BS9Ba9Z];,&gK0LQg=
1NR1&KX3g/LJg/EJNY)X1)0#AAF>CE#>V[L&4_DS1P56If4A[5AN#<g+1AOgE^9d
)I&.g81>R_ZB22,ag,=W=6VA=FGI+XXP6CcbW:=WYT&FU^)777Rd..??1Y0cfFeP
+SY3#VJ2I?K[-Z5@EAeOSD08Xe8GD&7LM.Lc[?9=g<-NRL^2VP69=+KJ?bUYH9J3
1B_MB1Mg1PDE4I4W/6,HSH.H9.WR0?OdT?]B/C<I_1H<S@^/We^P0;8_Y&A)[^)A
N/gX6@,>=f36A3?&V3DK71S)X[[WF\+]d#:Zf@fS:g]X_e<#])ANU#gR&[BZ6SO\
1+DJ#Z)/6CYIUJgV;7[\.SZ,H2K=HBF^()MF^I?D3<6G/dU][/Ha2TQ/=1LSaC;U
_C=6GR?[H3AL1Y,_KW/,J9b\aLbH^XM2U^/IV8+JM763d3&D1CL9(2_aD_0GW57#
>IA28YF@W<c+50H)g46:V8<V;^BS:ZA&+6,YgXTX32&,W)/WaBT/gJe8DMK7#aEN
b,=db,T+bg)DG)D9D\HO+1-/9E1QM=T^B)R]E4UM9AGYC(T27N58(?(:-[HT_^Z:
C>)5OM4AC#P5?2,PMDS:dd.T)NZT^aY\S=D)^5(=]9YUC3)NF_:=#+J4T,U_<dH/
#-8]S0>6(WDP7-=gDG6>=#0GK3CddC1J@K+MR/\T-AD]-@Dc4\-H:,3.)WSX9H2S
R3/[FMdHT#SRMVCMY?251F7;M71/9W:[JGXMfEGHI#fe>a)/fe3b=L[>RA:0>@7Y
OgB+&LG\G0/=IMA5&Y_G-9c:CJ#4XPe<Z#=gT3)BCAK9#Q2WAX;S5M6Z#BSR?+4-
A5#W#a#PeLA,L_H\3B9P)E?M.\DPM6VC-FLV8I@(:[XeL12^V_;eMZ5ED-OPTa?I
;G)PXYW?cB?Z[_[QSZVG7<c14=>>=GfZ](]>C\[^<+MYUI[(Yee]J]ACN2=S_D67
@\bV/4S.;71/aL41>#ADRP.[Q/9[GM>@)XccM98JKW7)CEXZecIX^)L?;/U4;NXI
]7f<4BaI/dL2?(@g/M2LTBTS>2Y9f=NXVS3dNUGg?G/e&\46,CG1Z0a@],20L?9/
YKB4<dbU7SIJV&FJ=e06/#94F;@I0N;#C()5K\5YK0:_g?02[/7PTFdE,:@fG[H6
>@;Y/MI_cg3+PD5H<)GL[eD9VM@3\g(J_IBK0Y3gJAa(<DW2J@Zc<TR1Y_CfR@.C
,_BKZCOLQ6\P.?4&_a3IGb;V#+U+3a_.gE<E77b.O1BJN\P5@#Nf->f0N_N,:Gb1
c)]HWdHT9/_.T:<Z)#Z3I<Rg/?0M/Cd^-[<4U<YW:J4]FFJS9WRGdJ\LJK05G6#+
PK@ZB#EJ&6A/;1d0U0dCVIUJ5SS(G3._X(DX-B._+:DM53bP:7If0^M3O5[f6/Cd
P=L;6N=H[[NaZ(e]@BG_#SJ\D+0);EXDL<EI2Ff5/e&>MAaCO+U8^BJ:Q_YN@?dc
MILX2^;VU)8;:c,-4D-O#([9PfV6)8&UO+PS\<aR(QV?\d(&O?a:58ECBe7R<Je/
b>CISE^P3A@_NK2S6NP/8^L+US@Q7cdI[+T8_eb=+CdX7O2.0BKb.&WPL^Cc9/;8
cWSbL8;W\#W87+IJJ=]a2[QV+dZ8D84QM\,f]KDE)GRTg(C1/E1(C/CgQ;ET<)&R
_2BAH.@3_P-Z_^&0)K.M(<_P2Z?=EV,@3H(L]]JEL5R93FEK>+_RaR,;JdZ-K.6\
JK>:47D(-Z;2-DZW2[AWE<5-McI8-IDQ@(49e(3aZ\C(bUFd=eW4A)\e6XI4D@L7
5#>b4^;K^<#EX6LLa<\deM;TF:dbQLQ1;KZUE09._;SG6g>,LRHPXHHRRT1Y_S^]
YR632-P8@M5EONXF9^9K\)(Y[a:=)@_<S3gQ?Nc<71:Z5D,_GcI8DJ2b^_GUUBYV
UHg6KSEa)cUa?G-Tf=U.\KZN,OJMAg4?/SN=Y42KQd2E65>FMbS/EWXD6UKM>T^>
[2aLBNDAUHg&[Re7cOO(ASd3Z?RTTOP0#A=B42-B+R1IQ#435@eJ+@E8Ie]HV?M:
U.B07EYQ5_>HIB2gNEMcV64[]]5C?9U:SP\3^K]bgeH@TZ#=Y(L1_9W]_#(1I;Rc
5e]G2E=6C2T+3Z;ac@@15@[d@N&H#TcD&TR2G(/LZLY2OaRZd\1cGN=0U)1V7^>c
-D9Q4[SJONY-UH0D^(MJB8H-dQW1]]GBD9-H53baBF.#>NUJT[GBNJ/T2,4J-NfP
_d:U46&O/<](_Ha4U&^B36+Ka063^-,7)PT;H8)C0ET]f9.17-F.H)-B\PNF/L#>
F=URTZ9F-[Y?XWA</VL7C:e>01SX^Sg<Uc1I>WQdTg(:Mg]RK9bE=<H\aeC</AUB
<.P0U;PIG2_=HS-Uc\ES-0?>2G(LKD<].>e.D=HT/Y#[MbeJBc0-7W6ZbCL31O\2
XJ)^X=@;?XYW&#.]9^3d.dH?9J4aX:d0M->1;L-.W[X4e=JeM;Z-&,R)L^7/^GTd
:CT<WXX8T>-ZKbg#bXZ?]GQ4-K=KI@JPH9Zf#;.)?K5RM0D13OM(Z(bGc,ZHQ#13
&R4),PG^+ET=2KBUZbC+DTAYHdMf(&(=Vf@ZOOJ_+c=M#AZ=0GRB;KeeQZ&g5.AF
HTdXd:-;:bcFPC,)_9K@2G:FB;0UaHDSgRfdd?:)e8WMbOH[a6e#E6(A)+M1C\\-
THZ#\XKCC=XIK@(G30&43H]d_a&fN(K6&+/8_GNH@6f+aW/A7+EaV=M4E\(DW\L+
f7@+(<8Kc-_?>R(;<K#OK#6<f>b@#Bc#[DJQLd^086@<KFPVV,R5ZLS/:OGX/7P3
D_\9SJDC6-W:ee-)d5cOaT#U\SJP7:f;+3^Xc8a0M_V)b+K7dPI>W&Z0)]#fP?\9
])_L_/@K?@dV06EM+>M/N@G2GS?XHefG]&FEM\c^Q0,0@OMFK_8I(F82^@Oa@=,3
Qf;3gX>5)7>2]C^L_,1Hgg[:8HRV,C@=TNV](CCSI.7]@Q3Q=93-FE\@Ke/Kd)(A
A-IIWJL.62eJ?GZZcOD?V[<WYa;#J^##J_Z(H@F&\M6c/L9OA0>QPWPf@=Q1D_;Q
_dd?QH8/W6BN/)76\-39de\CQ+9QO@bM([@fN&1cRG0W,O@S93Tb<9U7?X3CX#)V
NNZ8G#74aTE5]<_ZL>CAHa_P];A&-35[0&:(CIKY[[JF>HY,:PPH0/=O+6>@3E8E
B)c+YPBL.T&()5FS>2D2?(d+3e8X;e_BW+12L(S\aX<[G8ZNT<I&aZ_TAa#DJH5T
DA5.;QHV-#FLIX]b#WKBM2@-d7Z2+P?S74(Y:Z\VZX.2&(_&7_fO+@<C>4INK9gd
Z0+;6e,0,CeBG/0B797A6IS4H)YEe\V3-OR#YJ)g/YdW5>YNA>TbAEJ]@2C?+T7V
X42^f#cS#PI_b0PP+;.EaNSDRP+MNNf(V9&bPb905YX3Zb;agZc=7AS,3+\gC6cd
X9gg:&@;S\DJVDQ>Aa^&;GK0cI@9X30L/XK>#\\H5a@PfMB>(6+-G7ENVgD=VA0H
/RcHYIQP#/T#=7BMT6:G=7F,e?WC^0>7T97@9ZA285#6HNcgFTEO0)J6(V6Z>YQc
?T.&]6:_5I_G4()&bJNA@3/VcRE>AIO)X26JVPSEDFO57N&gO=Jg3d#N+NGC=U.5
;GBU\UX+J\&7UA\d:eN@M[bBce\FKNd.aPg[9gg?-PGE-ZCNY#>8e4gZ17XCN+V#
Q;R[<SZG,D#J9N[\Qc3DKHZU9WM(JJ=6?Ag0E7A0KA(?&^HQ8J-[&U:YAKZHFQ<>
#5IJ/.HP(),T^I=g,8ZL:YVCR[Zdbc1(Qb3LYH=2MXM#A&P#fI8W/#f/ccA=4(X2
YVK)gFC5)e,T?H(/fD[,3P+g<8F8Q6F28>B#784JB6QV7((CBe\+.a8#7B+BG9>/
@LLb9#L3b0NUbK;-TU5#((#OcTaeNNTRC]GTT>W<(d(:[__55719K(g8OOQ1>Rc[
A+&#KNgYfW64M;7d\H=cMe)D0@;CICY&-E@8XVT-MN4@2P2SQG,aSO>JI]?1YfM8
AQ&L5YU\3[\<A_GOZD]a+CC.HB:gYS9MS<;3dDK>ECe[\La0L9<09cNL55X0/)4]
+1Q0JW/YLA9]ade?#?:).IXHaJH=@aQc21)B;V0Bb8d5bF45QYGBbE;)Ze5M]/cO
cX2/C?fV^]VeAMY?Y&K/2f]H82+CL660#eR-dJLfR77TdXPS3R>,B=O7e61?\&J5
<S..[K&T9,bQ_Rcg<A:=-@ZC9YT<-2X;7-:EJM.)a;03P&9,LeI-\>G#2c#4+5K_
;57;c+(>4(VJ\Qd]4LQ;+ZV\75G5ERB;]HO..([4WV;(3F8d;RN3\Q;@JFda6?29
E:8\R-A[9:PTCEN\2R&)8&c3(Daa-]V7a5>8E+SVCKSZKU^<Q.,08=OZ<c+>PS^C
f#>TOD@ETbS/<6fHeFJ:1Y/3LE^9FMW7CeK8I=XR_P0;X=(U=&XT0SgP(C_F@GBY
G,_/-cD&#SI=\45N]-RVOYTFAZ,7b7Q-\L1AB,03gZZAK)Ic;a;2@-O-T0a-a-ea
NI5JS/TdHW??cF&^6OR1H+b5>Ba#,=R;P&P9Jg7RJ=M]Pc4NRY9:_C?+:@W0bA\5
7WE^59a\6,&eURfPS_eR6::TDJS>J((G+8\]GT<A#9;7PfS3eU[0#aDQ(]N9QEcA
XF8S@(.+NW^#UJW[\8,#Y[X-f,I#IE?>+=,<YS3Fb[,0PX=fJdSGTXU=,[QSZeQ+
c8&3<S?S/Dca+HYW+:13b1Z#D5&5A#O6?G^.5/J3V4KD-JW>JN9G],[3B(=K[VX9
_-_\<_Tfg;/(YIYY50HaSF)_PC]/WM1/3/SWUMGY-NT#<=13.<cZ5X2[.QK)cER1
;F6BT(#\;cCE+S3Y/SZ1=V:-WRM>V4)ZB,Df;4HBEXJ,+CL;<V5?P^,5PP4\^3FR
g8TcW>fNeG#+S,d;UJUNGUP-AKFSTLRWZAE213(OaHP>bTCATcgQ9Z:SG?4O]GC0
YVfe0FNKaN#e0E,T[B@b7_AF-M55](Q-d@A0SEZfHa\=M[ddSM;a>2d76a=c=Ic^
+K0Y?Q=K6TW[H(.AA9Z]=7Z^b]f@7[N>XIg(DU<ZeCe0ADYO55HeSE,d[:7Of,eF
-M-X?O7MFQ?4G+B@+W_HE(cABf5L1J9)(6QRT:7a1=c[Q0I/0fM,@_5Q0I-<-?HP
#]4[,83_fag.N1QPT(-O>8/<LDf.d8XFb0@U-BX1;H7LZJ2gJ)+=;[5M&P^6B1Z-
IC?AE-B6R5X4c(51_(Oa:XX54IH5UAJ9MP21,HSE,V^99@6(be^<VgVH&V]4Xc?P
>+V+Ec1OWKH>0N#9TRe268GVg\\O36Q6EDD5ecaTXEZ8<)ULPT[((C2TAKQC5-Re
KYg]5PRM3Z8PWYGTb=T.;:>\B11-6?8&1SY3WbeB2?dV-L0&A6-<930T)?#A?.]&
EaM;-S^(/I]KR,(Ofb-^S5JO,(I?HP:9ESfK&1H;7J1(1T=(FH+C\F5JW2TZLdN@
Zf@&G:^U-,-f?db9&BF1:=]Cf>>XA48AQg<OPGFRQ(-INfH=8@G+gCDMB)]aYSL9
CLC-eN8UCd>8<0gaF@TZ+138WO@J5;P@ZcBIRc0IDaW;9#/VS8N#J&-N1:4;J>&W
T;[I6+S^cP)f_[fd;2&bB4?26#d9@FG.7Va>G.8C7Z_1+eEW_O-O)UF<4TVbI++O
c)Y15_L[eK#/KQQ#35_e&^MJX#dae8=P0K7\C-,,eIaaDD[D2BVE7PGg#-HNI=<E
>b=b)Ig:[X3][?S@R,FgLWT8U1X/Vb#Y5V2XE5QLS5S;Hb^3_T@;HLKK_Gc941[>
9>03+9D/b2g4.8+9BSZ(:PdD&@C@e30b@Uda1M+5B.g@FdgUM=<@.:H?AK1_&#9-
NZ[Ie5S5P:?2I\)F_\J4U8SLdKDg/AA)Y=f_J8QS-FdEQ?.?&0#gPe4AAdg\>59)
\>77aX9(308-I;f8B,bf@bYOD4T,GVXYe>S=J,0=U]=CD9e5Ff((Ke2(+g)d7aVg
.bQS-[&</GF=(0A[+H<LV9_W8F:,288MK2F<WT0X1<]C/>BSLDB0_]Sg&^R8;.7:
J:(bQV<X^;BOMB_c@,2J-g-]fcA86MbXBB;GEMLW.PBf[VPc/,DF;a-3dg3?eA@4
P4R-#d8d9VX+=b>TLcPFQA(1g^MW[KLQ=#,c_#)\6S02FG)@7[M,a\c.?dL?AE0-
[Za<Pb1>LVM@>E++5(LEgB]1_,OW^UL^N;8J(5P;^PPC;9-e:.VK9D-JO/6]CRCT
Bd[9HN=XI2VJc92AMX#+G0U+]cAW[0+:(&-@Ta8ZPaD5Mb<8D,BU,08M3WF5\X?,
K>-ddS8[&>g=RL]#fgf/8P^5OTQc6a\PVFX?>H21?J?L#V5cYYKaJ8_+^-ZPa#Pg
6Fd@^cS7DfTP:N+=E8JPR_3LW0+:XQ7da&18M6NKS-/NX1XgG_>F=D0g4W.04#D@
dFd)7WXJV^?5V1JeWEW=__Z0<5Aa\e)aC9&Bb=EfH(_3-0fgGF,,<A,[EF^2Q6L0
G:3B^Q+@f>]7<-02VV)K.D\J[][9>b^2^XL#S[C.MA]f?>O[]1]de:NY4-e2Y6&R
;D2X.+f,9=L22d#)S_<1fV=0K](f2XHb6]dOE/cc_.K8Ag+SB[\<E/dG,+e/E20(
0;-c)O9cOeRW?PN#<9;O=W=d;QY9:)4Xe5^J2):9SER23R:3>TDA4dFM#;/&882P
AVdNTLHD\g-bWTMSWI/2N)c/f)g<7Lf_UYIX.56>ALA@&4fbNd:,8<=HT:;BFe82
:0<g5)U=^dKRV/7F_B@P^WZ[ZWIV&:I=?;GeLH[5AcQ2fU2=KKT#F)PRD6Ab2OS>
cR\.&,AIWA6(5B[Z8[-S=S+\#b4[/f@H88[45>6DLEMWDB[a/&e@TCUHA(E61fUO
5JS>1M9J6+d@A((?eH^1UN-:HdM+6/7gRR\VO0E,2#NQeA1/_bJS)Xe+L9RANVTD
S0AV[-JK[/CEYE)UW6M1#HEb[_,AGeMFF)]E?W6&<,Z:\G\G)T9TIbY]dLUC+6</
RR^1R5S0,\E<H8YPG?@ED.cWVCca?cG7=/SG/@2E-7^-L]UMV#Y0W27>(.ZWD9b6
X#K\N,[_X=[+CJ,52=2KTgQ+4M2M-GVZ@PRIPX3_]L,S-U(]:9dHcaMU:E33NR;g
D-P-Db=&2eT833A_&cU0),M;)@6N\E4Z5-Q0gF[bU_EM98Uf8bM]5,bEVPEHE)0G
VL.F3cA4P0T=.2I\>OZ-P7=_C,9+Ee,Nd-L]7bKd-QVU<V5Z)-cP.92HTBe201(D
+5NbH54L-5:I(V&6a=e<J-[dgN0B;GI6d#5&+)gJ=,f\&)6[WW)_H6OFE;\2a/^J
T7c/7X1O:f@&,GI?_;KfSX,7QbBS<-eO):2);9AW5M;/CP3fJB[[G+>=XEL380BU
3d7=XI/CWa0208MA/@cH0b4aAJF[f48LJ::L;>KJ:ZH4S(ea4MC9@/A.Y6@T#M<_
ZccG2N#\Nf+<OF->/Gc2O;Ve//ERB+bKJ=H5FS1aQ:a\/I3GV_/]Z#_cWdH^#;EN
TceA<\cL;-BA>,C4+<?DB:C7IC]Z1OP66JH]5AXP=VfY<(5A4.RYeCC5);6_,<MQ
OOSEG@M)J/a(OfgJ(?68Q>-g;+Q]UX@J@Jf(ZL.\((=GaTIa&B@)>L,7O@e1.B\X
H8ge67d?FF4FaH#.?Ue)bFZ4W/^;1)=Jd\K?cBEJgM#[O1>?XQR-24WHfBcb\FMX
YY]5&ZbFT2L)N<S9:86\I9;dE3F4@PSW^BNN7VO5>)M,5U2.:LFd95V_/.E#KBeA
IT#R_D+KH6KP5UKP;VS42B:(4ET;HXB79GGDK8K-1R)U;4UQLDY7Sa@AB10-)X,f
H/WGMCK4TS(Q+7MCa=c7R,_\;8X^]+C06N5.I+U[VMOa1A&1M?,g/&19XP.??=I#
++&aVf_-P@f\g,EUDW(&a/]C9b=;bTGCY@_OJJ=X_bQ,TRFAIDUY4-Y+IB4AGe[7
@>4(I5_+/?gS<+XQa8a]^#5W3O(Ybb)Nf9VJ<-A=2YZaBb/6FA:7\A;[1)98@Ae;
OYC,Z]9SQ@5J<34LSYNZ^AF^&1\IFF@8_c5E6O.;,_9gT;FC&/LMFKF:^10d#/9E
VT4VaTSRZHXUC.<::a@\EI;1QJ@H3X6ZWFWGHfO^A6K>?aDb3_U0>8OAGB1E=2#1
Q0:-)8,GF<FIS@R<7Wb?7U#<f]&+:GVL8+W<E8.YE(B#]fK)03[A\43@MQ.MXZR&
P.#I3UA&eHDAcGB3cTVLHU^.C^W9,2;(cfg])<T^;8@+N@CTb.AGc@3UE>42gccW
-L7SV<]XJIKPHNdS\#VgP[dRf:J4=^b92>ea[V44JJfA_BdDCf9(;/:<c-KVa>5N
:bJBX9=EZ6)^I[bN.-Ae:Y9.eDRHD):@AN?D_eXP-LS54IJ+N16)1c?8FW/eg?O?
MUVYZQ^<1)MKRN=LS+8_Q=V91Hc(188G^U-W1bPT)WC3^@cXO/0([&U64CAI2O_L
3LYZZaW?AZa1b,DGT#PF)gc]6\IBGDKaTVJ2F>&&/W^X.<TFUH<NZ_T;1-^;_:KJ
N\5c0cOGGSXOg-JG3<KB#aL\\,Be?#bVd;-O3Q)-:BT25P1fLT?3_Ed@-0]>Q<CF
R;B,\Q)N;F:BV5]2H+gOZUb+UM9VcBD-c;b0N\F\b?Q>a70^LJ82_]F5W=YUW>cU
6PDD2_bc@F_QQ27g)=;U&RB4F8BGM=FL@7(??V0K)75fV__?)@7I,a-5N_O3\@.@
g<RL@KH5Zc3P^LKI,_X2P.#P+YZ.Ad3FMA2+8-,E<\UbG=R?33-23BC[3HA0S35A
9<CY[&D,^H;);fMXbY\<WWeRC&0(#bTD92F8L#IFV.91GMQfRO(.-WLZ/-B+>E,b
KaMLOc9AF2c:]&eMURB<ccLT2T:T(T.EHD6CPYG?S9#+#(MVBI<DOZ;1MSG8]DND
\,^,f;JH)f@DQQ_;Hg.+3MU9UA=?5RgCMJN-0@>[YBebfO6cPg+1e\d[:#/WN0V@
W,f0GGOZH_V)X@TMPI=K=8c=LN>/15[:OU=II+g51)W\0N&B9RDAbS?<8[g;84YU
aWe4H#.^ZULNW0a;7PJf7(?UZHQSSS>(;Q?Z>Q[>\#LD(4#.;#.P=397?^E.<\][
)gV8&egd[A#64YTC.#5DaL\DT>cHeB1&>]/WgRg=_b@;#8b=Qg8L](G^;/Df]WC&
Pa9/D)KV_MVBMc7Se)0?)[Y\UR<@OZFU:ZINDSa\>=0HM1fVPcP[X[55->#N991U
eVWS.=8A[;UH1;ECe;^c^>U_9.b:3R6ecPFWa<Q8W&.bXgJ#L]_BfRM?9VQacBS.
CH@EA5>BM3W-_&[&R]c^5WESNB4J=K+YJa]W13>]@fc[7;AF)/QNE(T8A?M]2YYI
[;(@@?-FY68JRK:,OMZ^W#U909QRcGd_Y7aZBHW:S\VU[2AB^J,<_12[<,;K1M+K
CG]P3[V[KK+J@gXb3RfFHQO082TLZPcc),JJ,.Xe<2:P>V(H-?S58_0;N@,J&DPS
gM0XUd08:I.5<:I,Tg(bbP&=XB_QH)U,L8O#2I<M].O+W/A@#Q_GTDK)TZ/:G5ac
#5(?P[;KX[2PTc;-)U9KZ2M&3V,_P[R>+F^_<[3)>CIZ04Y@Vdb:c\[Kbc)NZ]J7
]gQ9W6;?eCR@Mc+@F1RG6/(8<Ka;NKDI\D2MQgBQIYJd9JG2QYX2UDTG1.A>d7<4
Vf2NSbD:gVT^20f:+<<cY+U,(U7/E1^-:ZH/Xg4+?1ROO5dUY^C<ND:(FbZ4;Z?#
Nf)V##?[\54\M](#YGE+a:@+.<U0A(4GC?X5da2b5_H5>3<CgP6WQ&WK7fbg&.GN
fR9C^V.MGOV?db)3<4=Db\[Y5b+&D><2_A+@\c;V;-QD[+&P8AYa#KP,(c>dO@2Q
;V94:_4VTIb:<<?&f^Ba6N^\=..&NV&<O=f13;Hb^A,&CPE=TIYaXOY/H+A+J?QJ
^e2[<ZKJBUc4PGD_=9_Mg\H#?](?/95=7I36(X8VOaW<0SA=fF+C/0+>C36]<N56
V+[LEe47.H43=;10\XSYB2QSNYB/8)W^gFD&M4@7X4.f1AG,OX8]2I=07OJ40+>G
MCR^YRbRII8-\R-M_,f]4JXW^[_NXIBJPXRE0]MKRe46C6E(WVP3f@:ZV?9G_+CZ
I>\F[T0-6+)A\#VR[c#D5ERE?DL\bKUCd9R3Z/0>e;TZ8M3#QE:)FXL#,_Z;MKTG
L8WC(.DcBdX:a\OU?MdL[87I.B6KO=H_I(A4+IB:_8,,WF/e6e-9-2BO6IU^\ccO
.-NTN.AeM21)K4dYf]K,MeA>P&EQ9]b.<M3L+54U_(5P88Z1<9P./+e;5?g6[XL9
d1Pg-2gfI\\[LXVDVWWa3X\)>+WBE;&RZ4,.SH7EGQOLHY@g-&GdX9CL5]A\3>3Q
UX#O@D+d7^Qc]&/BI-0M:KT93@Ieb9\BVYGP,=:K0W.gW:W(e4L-T?EUV^G#6TE]
VAH,H-5X@VIMH5Ve^?_BUVIW-AeaKB=d2ZCK3#55:P]T7SgRN=g0-[BfV#VEDX2G
:N;a06Y,/1R6fPJ,]S.?Wb=VJ7cX?bC8[W#:]F?<<N&4ZC,)eC8Q5A#Jc([[KbDS
QVUaFSc,M1-MV,Yg>:e&M#DD\U\Vb;).6R9U&__8OT=,AE@QQN3af0L]=e(O:GfF
\K=2NW>IITJB?DgfV>/SI:N)/]KN8UgE6=gcK_]U<O^>F5AF0;MMJcCJ_Y)DdFKN
&5HCCLJKLC1>EcaB>RY-fcBIe#f7#f/E(3)J=K--d>_Yd:H_+0O4N?^.=]S+;:P4
[<ZKDP/:J4AWLfTB>^+Yc#9HHV+@YH86XA9S0N9QULW)g_.=:)B.E4_+dO&_)7R-
_=XW=L\(&BU5THKe//@WK(3S?be>eQU#fR)XN4Y?1NQ144ME-MXGO&RZYOOBMf\X
=O4TeUY/N3.9@.LO)W@R.Ud^eg8YB9fO:3>YH8TX&SaI2BF/376IZ)c.+3YILEgG
X5>JGL1^\;10ASQ:/8cQ#V9IM6d)F]J0Fg]/\g<7L?(]/>H[Q,3FW8UP_/dLg<NV
T-aQ;cV2<[bDgP9;UW9F.H.BF1gSS][7[)^KZ:7e<7=9M@NBATdI81Q3K/YOSeD5
(P/D#<GVT?PZ571[9<)&+@8g2#E9UX+fW7ZLZLO>KS?JdSFYL^N]d#[I]gQDJe;R
-YO8ed,2,ZY1;;OObf@D2I20JZQKYW.<RU#.\Q=\gR2A33,f>ZfB]fX3JKaPJ]@&
fV.X/8-9Rf+I(O^T6PQD7Pfc4T#(.3K9[M0CR/A(O>g(65a[2dQ1M(PF(_EG;g+d
+W0c]<-0A/f.^#AXIGB+^&6E:Z]D7F1egS8gO#93e0#MU6.KLJ@&II)TO[V\01_(
R(05V1\Beb),VFZ0A>1L.PCQOII<>..;d]>0GV@M(Q)3MKJ]OLIUJKc;8^62F=W7
]CWg+LN+TT(&,.\d]0dbb)]0(L5_eC^g2VNaWa90UR.?c)0#0b]]>5NSGM9fE-eB
3\aY.GQ1&KL0b_,Ig<>.BO0;[TZcY5F\U5FLR_A<NP0Y,^N[QA#WZaHYBA6<a3_I
E7bT,HWGCD3;#T6=CE82IM-.D2\Y3X9CZNT[2I]M:c3BRWW;&]5_BAYVF+\3g/1H
]c2,fN]D>NAVLT2V;7fbXa3UC&+LZN0HL?R0H?a6Y^JV4G<#cgX7,2f:RXAKDARY
d&+M3^#Q8e(fRW/,[),&[[R_5aD.AMJ1gL,XO,eP;&Q_R;aDAbU,&JD&FXW-/f3_
5A?CaNd8RPfA73]ZWWJWC,2,E\?I>OO4<X>S<D6V+H)7NG(c[6HgSJ&DJaP/Z1;)
(Pd+I5<?d?U^gJc8C[P)HVYUPK\250)5NR8H]UPENZdH<@6Gd8H;6ZcWeMO4X,DL
4)OKWfD>4I;7K<,CM,0LW3dT0^8KD]1T-7MKQgd#dP9K&STfK/C)(6\AgTEAA/2I
Zg<=B,[]IZO1F[^E\3\Qc:4bMI8@=Q.5E;QL/7:8IdMCa+5ZS5163Y-aFK6I6]/[
Qf)b564b.X79;MKF2I]1CbHRQ(?7TX;F:.VC9&90BOPP8@95HHWFX5E,++gdNL+&
-++[,Sg^]_1P1c\4:_GP0c<;Ud)P^NEX0H>?2?5EK,cXbZb#f><c]dUS1D:ca1SO
OB-f6@+U3RCPYT->1bAM#U18);[#T0XMG?#XX.]FgP<2H/VAXRR3=E]7>8O;-).B
Bg]HH@7S_R0\X9]GZY6+F<&<B,]3H[,@XM89J4A.[&^6I#XZD2Z4N63X)R0gRcP<
EJCP;UD>W:(XG0WV)5[PS>PS-U70P_>L:BD.GCO]QC9Z1QYKV6bX3DAGeDWe?8&c
HPEL=O0:CAUaCC_:g/<:[#,ZXA7^H/CG9]?cNV[_dFRae?[08a:S6e1VFG9d^-/2
K?EK+(,&TO?GbW^[SI-YPPc)eN&f6=J6aC#8Y;,,O:O?bCSR;/e:@W\J741/7DH>
Z,YCdQ_GISJbH.72cI_HKJgLM=8.2EE#Fa-Z5?K=<-]T-<H3aAUH9;<MJUKd<DGK
Y]?FXBHBGKC-C<QGVIY.Rd?(KU^9F(G,H&egeZTEK;dfQC,9;1Hd#cT+VY?K03(,
?0;AWf1B[^e=:&VL:]PV)cW)KW]IO+/]VK/fPU-T96T8G&B8+#S>AYQ;M=[>GE_#
7NHI:3B9SQfXNC[_=XY,B#)gJF1?D_M\(GE&?G^:\X\H\X\OT(\6CX8SH7IA6.NG
COQ@gT:OfKQ/=79FFDSLC&XA6PK>c@?\8XA^f7JSPJUd;F.<C#O0))^eCWY/dU1<
C3T[2.7MfV5.a1bY3D7&A++0aX1VLNORR]MPFaJc2#D:b(0&:B^>CYD<,C,X?9LS
C8>-3cX#2&P(1\MR>Bf,XZ^6PE;PaCB;RQ1CVaSc<CS:_F#Scf9OOKBa<10?ZQ8a
9Zf4NO<b5.W@FV&0H^>NTa\DBFgW)6;;Y.H&SEM>/?EBXOG[H\f2fA[VMJ1Ia^+^
N._RYbI=,:@E3H,UfM#BFBWDe_&P6#5&W8-]TM&+U+ZMW4J5ORL634?P]P9M,)NW
_S_&D)3@-&bIO]b7fc@HcSN6#=6d@^UZfSHfOA;N&b\D\.)6&2M,Hd.YVF]1L\1Z
f+;3]<#+Z5ABBYe8:212[X=+W:DBJ+KW]e^.eJ=#Q2PMM[c7-X)a057WZ)@fP]41
Y8K84S^:IDL22gQG:Q-a)B+EK+YgV>R5PF2/J(D9fW#,<aA/U&c);4GP=7bA7+IG
FPQVHX]/)])R<+V[ILH/3dZMW?BP69+g7BMeHGfDcGENM[S-[E#>^4BXLMbL9H\d
0,E/Pd;=#S:5)9M)adP=\>F:K]EdAQ>fcgNB1Kb^eA)YcJ,XJ@.J6+TGL)>M[P7R
1D8@&;L?V.(D=M5H:g;6Ng^D4Q8=S9A5@,>Q&4eOC=L\LRPD]5/VZaYR6DU[^eNQ
RE]?U<5X[+6NZ2]9aO:<)gCVKfMEbKJZV8V(^U&QfGSP\Ndd6;2=KMD#7?R)6S&Z
)3P(YDbaX62RIgFGA)0UL.8I1f>5D\5VOR.=Ka5#PW#D84M5)/gOaPIADI8Xf)G,
3cAX.g+Y1.7<db@WeJD]XDJ;58:NG2A\MBOB9bHQ1.]5cPI>3</?D3CC92;QEX/V
H<Z5M>?@-b#<1;@^:#=aB1=fW4G>T5X[:d+5<(VSgS?-Z<KJM<0ZVN;RMQMDGPee
-.K==X/VfUI[E+JN##-S.G,GVdL;QB&a+S4^E.GYW0]VLUeNaS,d0ST:,_GZgDd+
:6IB7c#Y,WS^4+b,aNO/SO#+V/MZET#Y<&cT]L_747]EDF9R+/3(Q#1&Ce1VDd+C
[Z:V5)+GSgJX#/B\Rg.Zf5DX1a#;&=\Pd61CB[INQ:B8faJJbW:@B:>#JIT^11[e
O4AQcZ#O)NVQf627N[LJ+H8=D\^S3b1EOR,-dOGFSA7XM)(V4b&ZI?)7/P/5KBO1
UEIR+F[A[_g5LC5f&KVF<C4@C^26+.\-S[0@V_+G]QY=E#6XEbKR-T8N;0[>:O><
8W19NLQYWDZLd[b]-5\6U?IS55a3gRGPK7VR8C-XL?&PeKW3\b7#FXU(HbIdYSY3
#3GNc6FWcCJJ;FgPY:If2MJZD:9=_Qc^]g1TTg/=/5>DEQ,>_9c_Zc\:<76MT#8a
HdV[(_Be#M2H@Z\TL:2+DZOT@K,-8W=Q2C[d(KUGb^=a5J(cZ:RMK<@.@;9(5\#/
8MaPV:Q9AaW9#<:C8Z=80978d7_c55180Zc\Ad\]IE@&[[)A6,MBbL^?2cDX#I=V
W2D-GcT\4W^CeXP]?XOIZ-P/:fH^XA)WWSb8b5R<E(B\UH/gH+:(^?3HG?Lg?/44
A>f,(DG?OEfWcK1T,:KNf8YW[LgG;aQ5)OBK:8]g^V/F3LX748GM0^8++-d2J;3N
e=BYCBF3CU11MBF9]Q8aP2_E2&RS@KbCDU1I^>3MKV7fBOe2AAN8eW9O9G7ZJ31&
F(X[;WA5VM#9U2#Q;FB-KH@GVD-#@HOdaM4[DJXgEYeR[T&[HLc+Ba5L<KUf3@@J
L.F&#>5GN9^Z3[LCcOD6ULg6WCSLC:aJ_V/MH35I0@&]W4)>U>=[).O@#CM-0LFH
D(fTD:-fDdA9EZK[Ef9>=Bf[AY11E0CGY>g0:dI.f/Q,?R;aE>ePg8F;ISgY-?_I
+dH;8]XDVK(3ZeSJaURP;P7Pc-OV-c<^O<eec>feKM,cKbceeE53HSZ<NJYEJU=J
b_R1d]8B:Yc3LMU._?Cga9.:NcH@Kg4N70S[IZ5a>TNZUZ>T2K.Y_FaUO,(#&^.E
&+,:#<.c;ZKQ-=e\QWZH@&:C/,TWJG;FS:OSV=CXET;J\(;)ZP42\56&+P_^5bM)
-HGA71\O3AS]59;9BN=KP=^7eMO9fNd^\#FWMcY)fYCecX)(e/Se<T1FYf.U-RfW
e+&a)YG@.9+GB1[>:T;;T@K-T.#++TXRXWL.E)K7X4.39;;L_B+^+CGI(Gg6_T=B
#JR;4(,XW@HSP/-XW?ND5\V?)QD]M#@BZI]95aF8I5gG=_/RPS1)(+<\.&(J.f:>
,59H)NQ8Q1JNF=1GNXKW.F65eVN88NfMC7_IZWb6Ig.M97]^/Sb?V[F-].-17]W_
A##/ePcX[/.<?a@6aZQB[G@f4PeQMEYKaFf]C5g^:ZXI@Y.d2_TB\CUI6@K&gQ]H
aJOa3A,==BR+A\L#,<B4)JX&E;VMI0V1f&J&_IR-TA-2d7>QJIFR3\8^RG3d4];\
#V..:dZ@HTX)d9:66BHG-RM@_L5RJgb-dT?MIX>.^.a<aeF20^;IMf=130V2bU\g
7\TXU9/TG\gMadP^\39;O0_4b09>-C;>=bf;)L<\G=@F_?Q&MLNW>>#e5VV=.R_Y
ILf-g,-Y0KL)e<:b30#NefF-/@g8=^L1,T^K--:=LZI9-_9Gb4g:L=5JZ/8fC:@F
YeZbW\>/HOfLfKcY&Q3JPcaVLdY\QTS6>D/KU[#dA7cUcd,Ma]]C3_KX+NeNZBP6
W(TF\]5eP94KCX;)_XXKC=U-2RPKZQ]JC\Y.>28G5SN3[:?8;;gSd@dVKU@c)N_T
+KUag70IX:eG\A8JY(2HOd,(1P:GOF(M]1a/90aBcdC652gSbD]CZ[,WZ(&>=U/d
I#G@#ace+O523e-aOWRUI?-S-bC@WMUJgf/)&C0EMY08\DKHKQ69BCR+3Y=0:_[P
=WGb[P)DP_;7^;e])_AEA+U,ZEZ3\TZB2BO#cL_)HNVacGd8g5&;Vb>.G?0PVDSc
]LW@5#<#SbTWX[Y8Vcd),3@FE1f8M9a<R#-DPF5\P=<J>.#3fFM8DfW<-7=PcPF-
GCH?eRS(bW38A@;>=-V_T&DgJ&T#dE]UeaFE;,cF.+@+EL@Ia\<V49@=C/e3=F=^
=7D;b3[B=AMGeJ(C^#\UH0C2LU,L_ECU.b8C+G3/@2a@D91?JUBg?LAd7KVB9M<^
)[\&VMd1&M6T?W,DV,eV8c&DFbGA3SX:HRT#F6Yb8R-QP82J9W)A/C._LZ.L2S=,
^G2TIUP,PTZ&A+QGO&,X2F73/2=9ZIQTLDH@I=U-F5UX+;6&W1P41J1_g7&GRG4M
;B(](P:T71ba@eVKN;f(I#@:BZcZ]5:+0\(JAfDbcbU?dbBC2dEXM6T97YA]JbHe
W7XdC9+O^=:--cN1EfJ\>gX?J2V_HDQX6.f+K&BUb=NdbX>GD(8G#_7GD[Tf?_LU
=+aJ:]S,OW0_bdLE?<R[A=09^TLcf,7#-YAfFLe1>R@-Ce>Z2cU)[U9VME>]\(ZX
F6I#=(RJOS2a5/J>R,,]9XeLIHaE,4@HEPC;cM069aYT?\2&ESX2g2II,\d7=Rd8
S]f^P+K07MEeS08dLDf^T3QaPM4WDG<2c&M+4W^aKX=dZ8LBLDRcGT,EEEAJJ^0=
SD4AJJCS:G^J&Q._VfNYAU+\0Z:+-AUTMK8I7DR@[1c[DZO_LCB:)Rb/:U@3K<[&
OC-d7W#Z5PGgC9+>a-_#47/TJ0WM7>I46V,_(L4Z@.\A]NM\B\=8H_Qg-.6bgCHM
;>,E+cG<##eS)d_:(.Le_<,IcURGMdT+-)8(QF35+[_ec+3SO9PYX<_C>DdQ(=PY
ZU3,L5^G_V92E\+Y9O+P:=URCE-?^R+AGNQ0(8)T7F41/4gIg_Ped1-Ug[,C]#g9
_N(F(6F5]6<CYECQ])6P4fP\d>C+[KFbT-XA.C;JCRV]./I::a/Z_I5=O16B)C03
bF5TU#gT+4Y?#=edc)6CR^ZO-2.T9,SG?MI=HF[+_0S3\cM#?<93:6\FN/1NU,.R
]+,+<,?]B+#a^.aX,adC)/JAeCU75g])XT+e4#<B(Fg[=aEgN^J12dA]U.CU-fW@
)0E/ba(AT.&3;2A2^<:fJV=5Y@.KY^-dH=&A^-fgIdV6>VCaX,XH_)W5JCELAVaQ
UI@NR;K#KXf_.gY+KV]GLcG?3^fQ0R@Q-,^)ED8[BZ=FedH;?]K-SEGWRgDS?A\O
fU&U;?+(9ID:5]+K1:e;eBSf;PQ31B3D,)g,1MQIND,\86.EV[<f1&3=M#,#;I\^
@ZC<_V&0,?)C?;Q6-2C3dcA>IY#QbR&@dfbdJ:Z;Q=(KS-eJM<c6LcA=G@:PgD)J
]HB5AeWUYEKcP^3=B4_2#2UR/BFeeUc0&X\=L>RWM;7-8HKB8RgW^&0ECR=#00U6
+]XOe<-c#GXa3ZP8EdDA>d]ga:6)UQS?YQ[+YQY/e^bdaFZL.0<\I:5;XAeb2AN^
QT-6DJ#:1[dL3?e,^eH#-eb#1^:03^,.&b07U=><OC>=JJN&Q57\C,eC;3MKK+6-
=.f88Pd7?c;HeKM?M()(:EQBOb>?-,O[e07&T(cdeBX155S<,\33c_;5&7\bIKAE
=fO2_BN@gQ^,W:^+P7+Q1D&X-^I^fYW8BQW(S:C2A;YN>aE-0X,?+JSY&/^/6PE=
[_e(D\@d?:3JaJ>eQ)3T@P[393Z&0JHIZ_9-ZFcI&-e+cUT&FCeU-)]SU:4&dJ^2
.K,Q-S+(3XA\3a/(CdMg92GgY=VF1A[d+.YXS+0\V]VgU97d\/<ILO\5T;&a&&YU
d2UH(9JKHd@7]>Hb/@d1Z/58=bQ,Wfg(\^e2HUJ6<MB.=BMI0-82AY+Gg9-5(H9K
H>EU2eLMegU-:<[2fef@EZa.NTb(daa8J[@c[SBeJD5KP.2=ETAb=&0_J](H1QGg
B]H/J+Za];Nb@CU3H,AI,d^/)b3^??R;fgR.NQ:4D69[f5PHD4@dG=a.UA/H_AA.
c4bH?LQ);2f[XN2c]JK[X+5&U>Fe)?\UIWZ]?M_)g5AN[38EAG/N\M9&0,.^5CPc
g,&<6d]WX<FMOL4_-cSCZaRF2E)K(Y@IE:RLBPa<S0;HJGb<WW<ZC2>cUG^UbG;d
a?Gd6Lf4(RRcF?-:fF,N6BE:;Y8O?X@X39D?B7U<dMZb^&bUS)IIA,VND<cC,RE4
NdD;P-AIM:O);SL;G6G(;T776-Ta,W/\N-\0K25^,80G(e/g6N->0MAYBN#EZEP(
Ab;.dg8E2I:[7&>5.\IaUQ1MEZd/NU5[Y)ObOCL.]V92N2NB1fD_V=VXA2fD\+S<
Q&4[gL/6]CG/D1P@<MVQc+YUW5aFd&=F7)bD3\If-<ZJ9cg.&g_N:E=NPSf_b@=]
Tg>>U\;^8P,YVVe<[c^L2eKU[)GLfH@;R;I@\3BY0NJRR\^+BKH=RC_4YUMB2CaU
Z5YA7HT3X]+1VY-:VM;fIZ_[<;>KKYcF-7IL/fIXXWB^D@5\c6SI45@JWT]-6OEC
_?]aNa,D(TfFTCC6L[COS62\^IN.U7LWM)]Ng5a1g0@(E,2\[I/(AV6f_5#KLP6(
K:eT)#JC;II-6H8GGJQP;/.NDKZ,/<+/3BF4N#C1?B4Da3ZBB-M_I>GC5I:&U^Q1
J=GSIY9[g7\G0QZ)\^^?K7S>>QG:]Q2PX6PK-D>Nf:F_2CWBAPY7Fa8^1e:ZFcGQ
H\Z6Q3d4:WHNX+R7&R66XRV1D@P?J^\PaS3MWM5a2XX#\\<V)@eT_ULZ/B3fS\_\
BN?c<=SUKLUZKR;ULP9E=FR<9OGdCH\V85c#gEdZ_[aF#7?d/MLQ/)-beW2Y1?S8
fE+B_)=MTV@\J4WD?E\[U4ZfBa6+g@#eZ5fU??=5WI.7]AJXC<M;JU4dY?eENQRJ
W^a.VFN:&APe./a-/@8K3e;=,2:d#CcC6#J+fS/gFb5cVM>f6T)M+U@Ug>K&<PKR
GA8CPNA-R(C(R(R&P,[(@7a.Bf(C4Q.4[)/YD>be(Z:cRQd(eZFae]c<5T6aIK?A
1.]W?&C,8R;FIE:5(;(>XR+5AgT@7RUUO03?.NY?eH56<eDG(^Z+NP45RYX[(b2J
-b/I=;]_82PGe11X]@cBCW[NC,54<9;G=C^g+4=dRBK:@4NCN8JV^18>CHgGfWMJ
RRC>L&A3Q=05QMOd61>32.5B.K;07].WH1/N@16A\],?&DMMB\IE+E>OcN3S6K(.
;I-98f\1;[_G49ZY]Q?bDeBM&eE8V.7gJE47&+f0&R_D]Q]4^+;_-+QK?5CHJ:U-
,#eK:5\6N#?4J4>I&GAUSWQ:\PRHNA8e5(H?V9WG+UW?@>@5BcK#FVHAFB42aQ1^
CPEYLP9<ca6U;ffLO,XE5f&[V[_F+YVU(JZS7C#EKUYAP-S:_+1X)[Jb9YbaGIeB
YNU_QcP-&NSgaAJL\21?_/5GbK,35O&N-a,6YM2O#B9T/(:5)a]A_IGY\V6<KPbG
[,AR^SH^(2;O7(.DC[26M2B,/f5&ERYb=E]Fd?AW^U&K53/2H&N=LB@4Q,KLc[O@
G4,P32E2I9Z^HE02LM<872:7gea^8I&5YO1VU_+cN.X>S2a<=&[e)0ReXY+WQA]:
-EH)dDXcXRRL]HNZ&E[CNBNG8W.G<A28b_)=0^HE9Hg6Z/SO64\5+>&3YGHMA_f<
[Z=<c_@QWNZFP@8GVM#]DeG7DeDTKVaG_BAbIOSNKRD,GZJdE,YZ.dD7<;>U:c5V
T8c=?1YB,5P+NWA6[b<X.-R_?V:;J7JZFC.9fS?;@3,=YM:)a-4@=XZSNd\?<T:D
T<>04>.]gP7;e.[M1Xc8MSKBM\b^d5HWdKfTN+]8&2aF@DS1dKZUJ8(I)8EN_OJ5
:#CB]gO/Vf(@gMTBHX:K?[IS=F9HBXTdG9[B<\:([-A7NdS&D7/1E)H905Cb2(FO
f2eR(-Sb.VJT1&_N\P@E\dJNdb?#621-.9/9G_-;aFT81EJ.f&S>L#LZ+Zd;ATF9
[]P[>/d_ZWB9G?F75J.4g+,+Y(WTVD_L:S=PHN7d@c.C:2,;S?9LDgO]/J@DEDd<
bXLc5O/_<T?AT218&bDc]d2GB8J>W_E(AM;c,-7[0V4]DYe=:>1.a1Kd<EHd6^9G
M#G3WQ>)+BD:B)V/@@]9D)]52#:DNJGXc&G&Re8Vg2cQdI2P)dB1I#)ENQNUfU9;
LV]f?#^c@8+6AgJ?7((_23<f1,A0-KU(WbHKdUMX0.D)[#5ELf&PW/fb>EJfd;-4
\YJ[K=_9:-:[?daMDC]@,?1^(@:]P7/1,V:C0:-M3aIecOA7LSc<<(;+7T6MI,SM
:Q4Fg?e6\_0GX93N7C,4c[;4&M04+-97\8gFeK;17K7>674g>UbKg1Pe^gEP/WE,
J5_^N]LX@b&I(G_SS3&<H<Qfe5_Z0965QR55&Y@@X(NF3]eH-44<)Y3N^/;HfU#0
c7dEU)?f:]#@+dL7cg^\4?4fI/CUd_CY00DKVa/#\B2DBHLW]egH]0R;>T11)DKO
G\GGM),()Dc-C1SLHD6F94K.>WM(YGIReES#L_5]MB.-GeQ0?BZaDfM/ZdBSOLe0
USR(8[>adFU.e,W_AaS]5X&E,+,cE_Pd8L9f<@B3OZG0A&6)4M^.B4WCE8&P;6D;
A:Q?Cg]6Y)2bGRQcJX7E1LA9?/QffZ/gEVERZV2<U9W)e3).[,L:g9+7+QgcVbNQ
<>e9D-]^2<V:bMEYEBF/;-?Zf#45bD4Y\P6O+05JM^NQ#,N>?Wff;1>cfU4U]Cc<
B3PVH01LZE:9I29193M<;8[#<)QOK\A?W-KDIAK[MR@V.&_,,LW;)2>a-W[)-66>
0<FeIMcgD]YJ75A2X3gR=XHa@.6J<??f[aAG,8ZIERC^e]WRO<Y1@f)J;_X[FCbC
A)fM/IM1Za3DMZ4+R2@5GI.]/<X,4ELF#VXbbD\244;^H6:I#H-GE[4H:&OZLGc[
)U=a93-FE@=KQe[/=g[LK#6N6SYV_7#W97..QES+QK5@0GQO6TI3Za\ZO90PA-?M
H\WS&P:UUI-fXZE#GM:D<f<S7fG4E@53+IXBMT-4X^aaY&4&A-WBe-a,gPCaUW65
CSQB1;AQO=KdCLV,?De0S+O&_3B73_26a[6^Wa2dZ-G,EJC_EN.Q5G]_JcEb.>F0
:[QBD[WWAX]e/(M;3Y1edR[_/+P=/feIF48Z_TefN[b<fI+;@LB<E^7AA,e-Ve^)
<_SgR42GA]#CX2/L/5UF@B2W@4@^=D>_\JE7aSV=+@^VV;2)<C?23Q:_E:>1KeS?
cOZCB,.8BGSE+&2]8QD??3,8G]AeQ2[1>Q#dQ7WT33XM)^c>L(O.DJ2#4]9>XX\4
fE=8fdg<R<a87+db?cU3U:+EeB=?a,d,ND>:5<E^F_>PP252AD?a=8\Y#gB[bK8d
E-_W&8)X5bcI/AKLWD8bLU\,f/bED&:S)&bR(feR:U8-^3AM4,f1-aK4S#^9K9-&
EQEEaTSaM^P\)eP95N.5:fUA1U94Z;D,fB6I/;c.&&6=>3HcQaUd@J5H9(O_I8)X
AUeZBgg?,]dEdKb&AT&EIWMSa6E-W578Z8b=+Q;MV&e=aU^cb?YH0f_U++K71W_#
+_d9:6LMbK-fPNPUe#VO=+=]cd]N0J^VGIg?g538(S0B?QK&5FPOG99#F0X/c1MM
0a)M<34eF[(G:<_])F]L>UVPP)+@C2eP)QV:\^KBJ\d82-:/KLb(AW8(U\QTXTUY
YI8/PfK2E6G5)F0B.c4+a^[Ze6W@fJ^E<DX0aI=PT@1RG.M@9Va6?3/T?JKRRVF(
CV3;KB^>=Q.9O+FQ[.K>a+0G:Z:87QT4S0DZ17P<3(IA^gA9<B+&[ZFa0Gb\L.#d
=7[_YV8=@7[f\25/;4/<JS_9FV93+)f+50ZP-SAW6bMb9]gM6-4bN),B&CfWIc71
C=eAZCgFJXQTFDEDZ7/<LcXa=V+dZ57.(D,VPd+2\=\^HB);P<T4Yd9E(a@R=B3R
1=6HB6aT1&>,CE9^A87)\2[L6Oc@S_bODUY^>F.:(#456+1HWRVg96M(7WP\MAbC
D5>#7e@SK>Z9PNPZ,XO@4/a>89K#Vc;9TX/#8.8g\fTO8B]@a][>@4:?;2MfAU2,
<X9GD(.HR(/AU8O)_-A[eAK<M.@70;>R]&>\=#<XYW?5?_&?e2<XB35EIBG]8bS=
/_CK3B#HX]JO-.V)AF(W1<[R+,/aWO7G],/Ie:X.cea_L(YcT(LQfL[6&=T0^Xa<
YB.G3<UfHeGfEN88NfNC\EAGU6gQec-a(6^[D6A&DE]DEJb#)M\/.>)],Z(PI_B=
ZP[8GK)8NBbK/<?2751,JWW0/6CG\bOU@:VWL&.:gbcM59Q]<cH>gH;D_;S;6-VN
,=MXUIY95&Y.04d=SHCT@<eZ9f>U6-TdN27JEVGF69-DU:2d51SEgHPWO_X#W+C[
G00Ida(.D;eVH=,N_RB#FIS?<C8b8O^Ba)P<Y2?K[OD:EV2XZG#/1Y7X)4E>9/RO
Qb:GAd0.G/(QMSPEeZ#A430)Q(@fPDV4C_,:24)Z^.<L-TdB.DZ)4gAU4I)-]J5L
,/;49ba[]<S&[MXRXEU3B8a^Z&da5/P]),b;Y(4CeD[]A:STJ[fB]]U:QG3F>A8>
5XJbWc/9(@c\X//bUN1]RMHce+4Edc+]G\DQ5-=/OV90D3L4+SKfQg^c.G#g<;[:
cT#20)._5G6\7/>C:ZgQbNJDR2N-_U&KC&N7;E7G9e#2La;KU,+C>IA[0E)SUAXa
=:=M<IWc&S=f5/U;QfU/VE.#D5dLB+.M4N-O?V5,\S8GD^f4&CMGJC+JM:;E(9=;
QO^[RU#L3?8P@(+AI7\3AO:R;LV63eNYJPd4>CM<7X,DVPPPE&MD@]Lb/CNM\R)D
_355>^;YSQ:\FeeJESDPED&_DdC((H7M9g]JdG(Z@X0,f;SD2H.UF13N-X[f]ICb
1@0d]PRbYVDJTK>(B0F474B#D=L,eCN8=ETM1)G+71R4:JU00;^);^3RR_TbVHWB
L]#e;<<9?CGQ.aH4I3^A.6XDgAB1be7-g2KQH=;A7)@CcRH9J2bHDY#bge[e/58W
P)_Z(^ad#7,#BS1g^E.314R0Kb9cDYAP_HHb5PVDYCRT6BDJ6\Gd/bKBe1gMgBS>
2IGX2V?4MZfGK^VZD?1>^^GQ;D9.eSKVdPPG:<O.JXUc&TU(5W+L)NLWIE)a^1CN
^4UT;#:A_#,XJK(M0DTX9M=bF.H]4GUcb@\(=@5=R0\J^^OX8FPc>cb=L>=9H<<=
/Q=RF+-DcCW/U7PBW/^=U<.]+5U_aWE3[34KYdGRP6QeJ;?97XW05H5(O#4(#a->
+W?&?,,8CZ<Af^^/J1](Pg_cXVD;@-(<\M9(/5D4Y6HNQVEL8/[U^:YM[?&CD&S8
M0?>#W_d#MLE.g?;<@PL?Z5AH&dZ\A<LF(FQ^O<=_eRa\_g,\:UVAJKf=_Nf=0H&
SR9<5RP182_#3B^a<-.?c-^=4^A_R[2=<3_0F60WS:gTYFN#NHYG\Z9L_gU&0N;C
G1@Y<Nab):]Y5\AD-0@b-.N2b_S3cce;dSXdgV-ISD/AG=/VZ\2+fS^NY/KDAC_G
RA6-_1=<,7AB28V-U1^(RAPSGS4),46TcDeZO+?I46A\5>?#]F4NWNPK9<B8HC40
3V3g:@4fG\,,,8^.60\H,=3[)B=X>>eQX9G_&eEJ-Wc]]X1d6N=<Tfa&D>4_X@6^
&WM88\<gX^>.J]\&bBG.UXIY76SHPgQ51](JaX/06Q0B_>9Ocd7b?KNK10G#J39D
+I(dZ;[I,.+W3Rec(RfO(F0c.6HJ&B^7(f89d-AU3Jb?,?^4d1Oa::T]&SLLL]B4
5CeAT/\VC]0GCQO^JE_2(KUVK1.CEJR[CGNVLUf2Y=?6dZ,VGC6+YQZaUHZ)V21W
U/9AF<2=6<a]_&SL4^?Y#0//g>M9PZ-Y<EI&@PPcNfJH?^+_+C1/DcZ7_??1IU)Y
KYVD/b^09e<&JPEGO4>GKd6N(cOM29)+aD)R;(ZA)5L(>B?]1H;5MZ>>]#,D#HgQ
DHd1\C5RA+c.16FfAaJI[H0M=M>Id1ab1HXD&PgFR7ga.UI?3SfRB+)Y(./Z)N0Y
^]FJK/489/VJKD=4b5Y,0JHY8]@c9>cE+b)4MX56LUZB+_\M>2Zb?][T3/d_JS46
=+K\)^FX/_e6SN,_Ie&8NWXbTM3\/+XV0N-HI9=7NNK?bY.Ab-NV98dS[:FT)GB#
d=?^2Q/MGE7_IPe.)L-;AM\ID#fR,SAAZT@V,gdT:)S<=LR6C>g3E9gZS9#T(YEf
(ZdZ^BY/)gU9_4+-e1;>GPA:H(#HgO&JL)G^G6)IU6/.8BMeWW,+-)+[bF?.RM5P
5I;SB]CL0Z#6&DEP-;5Jc.1&QS;8@GB&RT_IU<EUY_;bDbI+2YDL@M/3OT=Q3R(I
.1>8GLL7X1.Fg=0_1#M?VI-^?;cMD/Ee/+8aV#g#Ke0FX7eYbP>EIX^^9LR[7^/L
-[a6a-ab3V=R^R@K(,Q.[X?3Ua41=DB@g\5G(AZZgZgf,.L,E<I[8g,@\f=f3#gI
a7]g0]BRZ5PN43D,f3U2+AZ;=F)Xb2ZSV=)9L9a1&SC.^?]ZTa6-SIb6:R.e;N.G
E(c;7]<Dd_U(Ed5N,RbF=_]97BHT@eH;4R670WA0O>^-S7;I(YS0:6W^F5KSX1QB
X#ag56DGLOd\Jee[E)GM0K(@]E@+2)3eC]1:B=ZG#7:T\/Ia[fTCQ=KAG4=7;=5T
H2Z#GEf6@0[IM\6Z0BRLYV(R.-\?\79<,4XFJ=8aQ]8R;.\D0V<Q/f?A,dg4:&,>
_JUJe7[8T/egcFTIeTUX3QMGJ-[H=bPYIE2HK^@<(1>^OP<&cBXSETg8O,)YOEG>
VL&HaUDL7aLH0KU?#&F@)[V&7WHaEH.[SNYJ/(/Sc<)36eO+91MD/?6>QL&fe[2-
./b3H1J)4HM&4&4)WQ_QG.BJQD>LPY6E=P/@).^5SgSeJYT(9A+W^dT?2][gC)e>
+O3_+2K]G.<aWb.R3.+RFEOVg/AS_g&^;.E[aF(-fUC4<?-/-RX4c/Ae_JOVXRO8
/5<bT5JMLFfN2IC1)873212e5&#,/>>4[.=4-?-Lg;bDYfaHXK0S]4R;9E2a7YVY
^9RBTId-dD&76WPD+EKDeQ^?4&F1(ADJGPc.Yf\c-Z0ZIC&d.]UM\;=T_eNRSO^[
@+06b9PM(.PV_4HEedbY2U-8<C+W5N=?U7]@C94-F(^TSO+5+5g8f+B7eX9/\0.\
\=CEH8O1HIR)A[:Y\cY(SD)E2[1<R6]#-ZJ3(3>#Gc8S=bO:.AFEAE:[+fI4OYWZ
?cWU.15-259EW-:<f-a8O7RT6QRDAD.(#7G&;dba-_>09D]X1[^VU,UAeT@9W6,Q
33R@[B8_bW;8B^3[EK)#=BM/f,a>9\25&FfFKB-]c3YD]M3X9I>a>=BR0P+R=1:_
+J26WZIQ.JXINe,1&9/a23J_OG75;;#<R=T8VI=.#-\D1?:>)7JOeFK,a@HX(B+F
NEMIFM72>@11,J9UQ.cB36RY[H77V4e3<6TcA]/:UdZPM^Ld0Wa@9Ya+:\6VU35T
)26]#IO,a8NVCG)=)FTb>Ndf5K)K#_LfL>JeW,Q+6D8DI:Mf6QeEcVW]8>1:7dC^
?0?U4R_US8>[4:^dfQ_ZIFZY:Y6L#P0OV#QAL<8J([_b;d:^R8H];I>X_aa[46_g
^dLD_4BaKYEa\IWL6ZQb\+J/P]4YUeOLP>0B9cT3X>e;GVPYe/9-0J\^d&P&^<N1
]R+Oc\<ddP0FIeI;&a2QOS6\DDfH0K7@)?g9+TWRP0Qa-S_NHAP(Ue]<8&)[c_=/
Y=WCST:\X@>3(@LH7ISdEE1)2EPc&9:E0T7\NMCQ8PdfKL8^LH.2+QMdG8\BU+]a
#1K=de;=5e;\e,f5&e=gRFE0R<;YE>_XI?0P0<ZcQA&.gYC4-C4&:89\)3\>=fTA
H4M_5MBOZ=fA,3fH<L)RZ/;N:PSQ,W=;5Q_2KCUOLI]#)7ZE0Jf9./3^4L--D,D_
fMg4gHM<(-6[B.H[86+]R/X8d,UAFVfF9_T?W#=,L=2,UbWKeG<HcES1bc6QK^],
.\O#9NGK,)3@NYLXD3\Re9N>,5RI2QgENIC3AOSfcGBKJ-?dfT8Wd#Ue)cZX7H4U
&bP=J]N[NI/65-[W381CaRM6W7V4P(RR?:ABCNR],PA>R\55<64/V4<JWU#F:U<C
,\YV<;T(@-K_cA]-gdD4e#UT>]MVX-PdU]W)_\3+?ce^8@)-SNZ[4.5Mc8GA#KI9
^HZ2\c_(J;A0&A=(G)1ZaB55E,ONGD>:DLg]9HK\C0J(\MB3MEFGf[0B?.IC2bU]
F:0JU]<a9aEBbU<OJEX2g#D6T8D[X0^P;Ka):/OJF>bYL60g57ZP)Q=3=1QBE_T]
g?bg<(CdefJ?M-62&8]3X)faSYE\HTZ;>SRIVbN3LVX@#J)[f3+//5)29>^3Z(YH
CS2b#E6_7?P29Z=IK]K@?_5+e<H/dH&^NQZ(RP<+XKd6Fa1L>f_9)&W8F8>QdcfN
.(>(:_af[7CcUOJ]47aKYAGTX5MM+a63A@9/BGY6:MPX@9H8AJQM;::QS,X4gG,W
;SM692b]L6Baea0c\,EJ3FW_I>I7O,_@H^_;4&?I[^W,?D7cA8+@/<=-SK;GWC8+
PCg9=.=BgebB5Wf(^cAP@LS#=\_D5.[8OZ)2RC#Z_EVfS)^.XB7KcTHBJG]J54/C
FPJB[IJ06e74??4FOV@aASE,WI;YV-P#C^YN6GXER&22OEAP(MeaId:/W>dRKLDW
,2M=Z<;bD][>91JUA^HALc<Gf0A_7D.cZ]MV<9LeB2a<bXLOEN>b[L]EVXT@_UT1
7ZNRbfCA/[J:W_b#EN(7(.d;SY[XfD9_Rg.3D7D)bH;<C\Macee7_X^/e]aAU9:<
M6[?QAT:E65aQQ_ZETE6C[C-[@-?2RR&SC:c=6fA\Ha2bR_>TVWS#4/@:M+&4E1[
6TS2+60LXC=g8e:<26T=G+0(HR7F#7DAMP,f)?C9R,dV[)@g(N0)]3+9PTK-;gTB
Ng12cbB)?-3c\LD1L(.AP^a<bJG\Cg27]HGX&/AT<OQC@-J<._.e.7FT&b7:M25E
L@V#bSb:N>3H^V>gH59+4;JF&NDRL6U.b21654<,X^3LHCT@-&8991IMd&;JVOTD
XG&LG5N@H#K2c&C-#8a4#.4[32(WHeDPP#O-U(7D:V<.7Nce0LS;.>(ICG],RJRU
4K>^.-6ZZDRW<c13W;CbcU4fXIL<JGQ3&>L2R=&OZ1[8]B(9,dYJ29_QWJ0fVeC/
+>B]S@^;bf&U+g.TfW&=JIH#-Q_d.><J8L\KAHeKP610SIb?e#/,58#_&9IT&e>-
4#RZH-(1RJ]W6@OIK.9?=?3#^S>OBY9bW>&Q(T#9b@:Bc]^Va1EafUA8+VIc\8S=
g)2Ge4(E8:1Z4\[P\YX=YE@;\1WK7U)c/D,7S2aIe[1+Qb_\[@N\;(?g/f\\eGFZ
\+PCPCG4-8N[-gD.H-\.beBG6\Z^Q[@G[CCRS8?N?:WZ\=ZHSc\CNOd>BV&0G1B#
g,>R3K-H8X(GB]f4;O^(,fcONX_L#,.N09aA7f#JXE@03@J&K0_\_NM(N,,HX=3T
b\90N[+1]dB9/DP9F[,\Ma@c05NdKN?+E(7b>?4;FNG.2XJHD4?TT?LXH7NSK7cX
GZ-LdAZVKPXJ6Kc+1RD3K4>A@L2:HP<TgAU#119WFAY46[/RdCKOKQ647J@>G)H7
265ECBBIOM[P,[]H>b\NWQN;1SEe>.^:bCW;+?1K@,RbMeWMG2ES-GbC+YAW>Gc8
M[X21eIFBW=A^KVaTJ+JgTG\(b@\1=WJ><^+&\WE6;(Z31:\JZ2@X;Lba,aZ,Y_#
P+99<Yc>HE+^#C+;C^MXfTcF7^_c3=-\00bGUB3LUW3Zf&/S\_/C9;)K>0+DXVXe
AZfEO>M1(d9Da?2DX.f(?(W-4P84-WP;2,6L].47@;#T\C61JP,?B6.-E/1eHCUK
fSOcER7fG0FG-dG(5CSV,ZPJ:^>^2Se<A,bA_?A\X>+2?@FBFg[M,XJ(<W&Y]=Ff
1EL8Hc[7V-\HND3AWbC:O1Y8LR+=2306&1=<@Gg#T.0/@XcZU_E=&4e\N#XHR-<g
bT6REa^\9c_3b+@K_JJdM@K(1.PT[0UH@^ed3]N@5_CF-/2)g_@^]:3-:O[I_P1N
MC?8B_-79Y(\g4WS\^Nc3[)A/98=].5;Sa59dcL@BXD?DN7dD:bL+-_CBWU=1D5<
B6E-1K]1[#D,aP9M#SQ(N7KWf\X>Cg7I8<:7N#6:R/D=)<J:?GRR-8?5ZNfb?T/f
2\C@]:0JI>>\b=ISU^;AgaO,&PCPdS2;VBHDeQ)OUVW7>^MMQRG0g91+a0/9@TE3
=WXSKgb1(.JW?D7[4W2.X:TJ3H3KD&AeILe-bT][fIWQbLH>1-=/)TZ5L6\I,PfY
<G6c-ea]L8@a[?M3_N6>c@.2U<F.JY^_G9HX+07R]N+78-d+4da/CY2P<9MC9\gG
:+?=[?gA#?MIA[K+U-))N3^\^0;FTGK41Y#Re1N07(<9(^UOMFP[cJ3=]/MV4WI<
d_#1\<(Nd)SMA-c5Vd0K5.S#5(c0FX,69ZbS6<C]15OX4@4_B6@dG94<_#_VHOJQ
Y&63f0\_ZEQfH-LNbD=d;6M/JJL:O<I+1c:?IPU;3g<C)^&HXXBZYEO=9^J1PNBK
B5Hd:>c[4dJY2ATb(RWGZ[2J@Gg(L[?8HaKZ0WMOZR\W1#\6@R9ZH=-SCIKV(.bK
3>T_>XSX[:+.E4?M(,X.]_/C_42\WDbYb8JfYB1)<P>TFYIP3FI>VPX8b=2U@Y[6
8]MMQf9G&A1KGO4.2?@?J;LKS)_a#Sfg?OK69Y.PbMV4,V4?4SW]L;Z;&HPAV0&4
1G(IFCYdE(QbQA3TcLc,Jbaf+4RM?Ce?M;1/=DV]af]586_dSZUXGB\OIE;HQS7O
#+UCMffH;D2,UPf?4;3eaCBQ\4\O;IY;K)WR(MJ71]>C2&UXKF#Cbcd]DM.P]fc(
6COMF7FfHgI9(FK/VAcX2c,]4d(@JK<N_fNNXT(ED,f8;</SBX=&A)_GLaZE<4M[
I;V89T5Y)D:d4CM&&O)?0Y)].[IC>M_UDD89/NfV]F@ILT_)]YB<_Yb\.e>+LPTI
.g36@+D+J2(VV4JFIUUd0.LND8.+cTYU>N9OgP?1H82#5?#=O-X9SVeg24F(#cLF
A3e7O_PUG-H5QK[VRdSTKbMN=7gWHVHGCVgWR0C9NKQ[bDJ18Cf\W:SJN/GC^@+M
cf<-(=[9.950@;e4+-[g\IGO6HE0W=C_G>T@He\[\8E6VOP\?G[_fMHM)C/PT?);
Q3=J:I#Uc_X+C+HJOA7&ePZfd(bLQL&&ZSH-A:I6-3.\&:d-9Z#?N_1g^KM;.9^:
cII-]U#@9NF8WNS##YN36ca>gO/#YfT<:AFM5faM]4T8M2W4-4212\F>He5RI?DG
)H9/P0=^deX;M#882/\,0#F>4c#;7eWc#0K.VG34C;GAF7RUN;\KC4Q#B?JY<KU+
;E2dC@3I_SbHEd(,_Ve@HG#]-cd]L#2b+55;HW/.BV2,Y\90]9QZc2NU]WO[=gEg
,591WZ?#Z0\OBb;UAJRWUGd\YBeG^cgWB>d2E_1W8D[KQ-=V[PegRTA<&?DgH98P
fUgALJgD9;14.&aS,&7?b/24Z.G?W@&3_[17?cLA#^HAY-S:,=KF-6),UYJO\?=A
2KK\H./[/&Vf+XWRfRF,L@N,b_:?,bZ@#[=/;-IU50-95XT>_8.?@B=Ka/Jd\5U,
<Z:UfB2XTeeBCe.OD(_d\[J5_EaK\E;A0TOAXW;g;NfXV07?:><TE@eCRW1+LG\)
>24ERYN^aa@^TMVC/fK\744_S4EM2@dA&KLfF]TRa38UG]Z;6I2/EHH;H8GNCY;W
9dA=T:fNNGB=fW08QQ9d)#;C3-79E.?738H=bT>eT5#A7;+OY>Mf61,/TS0&KWYG
aeYM^KfaF?.#C619K9QKEZ72U#aa;HVL=FEMCU<2UT\b_R@<>HYaTHRWK8aceW=\
ba:5DS&c3M]P?(U9@bL52^dGHJe<[H3)VU/\M=(F;b=IMJ_IX<3S98a)OfL-#VJU
23]@bIfVf;e;VR;4.@Ua[(UK&E=HfC1DR1].6VO[Y(Te(Ea57IVO377DK<+.#(8@
#0F8d:3@LeIB/+,6NaJ47<YB\)Ka/GWKYN]/d.-?cZ)0:@O4]<H.JbN4[;I&aP++
K@?Pb#(Z?6J_]CXcC>7>TMIW:.FbQ3T8b85LeTR17G]DP-Qeb_1.0c(X\WQO(1WV
)YMH<].T+HT2H[f#:/]8ZT@U2G5KG9CfE<7#dBF]O7+e<720)D6[J]G..QgE:XM)
f;A?6I3Q)KU12D]]U1MLMQSfW2S8P3BfUE3Z>J>D+H2Xd@edCPd^?XTS&bIFA/-X
WGZRF6ZeCLL^/0?[W=MgdDZ7f1)(8bIT6:.ZP?VPL7g^40ddV)gV7>G[;=eDZgTd
HEZ&?5(,aSQN91N27AU;TGOB/(/GL>1<dR+[<9@VYJ).Y9D]b0cfXDSO>^,+ETK3
(8d?.EF:e-;@Q_&fLG2LT>QJGG2@?d,=E3\MAa1AN9T)6XJ:eN/Xg#?8e\97.f\#
8@AD]/SI//-DW5S<+4;QV6-W@]./XAZ#=P5:HRSDaHKHaM3Q)VL[ZW]^J(99-PSU
:Q9_#=)HT)IZ_N0=a6;7SBagM3d>SG[8IgKe\)Y/gV92ZQ+9>dABb\fN(<(M2Cbg
cXMPW?+\@:^R>]R]<J)/A8a3ae>Tf?=LP-4B(WDLP;8CPfe<:J.B;XMX];?H0U1[
8N5<HIcgGc-O4ZaQ3?P/^()U62Af-))XJQ/8K:QLMHS\;JW9=OO57Gb]W7gANN-R
gdSc.2&=CCM70E8;)+>FH6L3G_(g<M0AYGC>>,P@<G2_#&4CS5PQ7g8.^(@^6@ZO
>e0W_Uf^BM&7DV7Yd/:We7X,)>KHU,5Xg+R>U5-bfF)A0[?#D88fd=53/8+@aaJR
)Ab\=9T?]XYccSQWQMCI6WH;@-G4TSU/K8(X,>Nc=DH9e\#dgN7KK\UDN7/B;c,^
E>FfGCVa+@]2fG5MAaYT#,BKW@\YeTe@&8W_1cd31HZYSMIS1@R_^43XaLR4aH3Q
]cGTG=8g:(=):14Z[#6)GK0W,?E(f>DK0+<<Xa&N7D827ZU/TDb9Yc?]6P,D^)OA
TH@aDCYM[9.VF>?JR()[^>:b;8E-SAU1f2E&W[+[g4-L]CNQN:[a)f/ZR=@f9>6Z
#NWIF)R)ZHQ-S9\+718=F-g[1\1X9ce3f6_IKW279X@<F\C^J>)F<cS,7J3J\P[G
R\Z/I)R,a6M4Q.=(_S:PV(Va:>GR&/CZ?GAPMUJ[^1L.T,6e\6VcGC1W3@X?O8F>
K\@c&]fK0[)3#aIR##51Q?0^KV_,]-EQ=XgU/ZW./XgQ,K),=J8K-8A8fJQ&0/_L
+--EHLg[<2E;f2H[VKFWBJ/^fTB]TDI,<R8QP+V23YRf3<<d?OJ(ZN\L/UU[9E98
\F<Oa#QA]\/HbPNTJ+H_)+OLQ<bJN=\F;W4BNcbc\^[QKN_PXY.bDP<#[cOEY\g4
]DTXC.8DT[F9:,\3Z.J]>f2R[g_CDLARH<cf]]S)H1YXbVDIf1dQY#gd(92eMUe^
D2c?3dBIEKA73#:?/9?STbW+.<a=(2cI3^HQ,#M/X2066<#G1-)-:1#,])gLH=D]
.VT><MZL=;8AGZVP#6?<If=5DdDKZP@V1B:e<6ZaN)aLg?-LYggW[@E>7g8H_fNB
F]KYa&49\eJ0@DYa;/&[O)W-f6F)MX23)M=1?gTJ?5Y2;G9>Td_YUfBBEX-d34][
RAHK2#c@IHa1;>:FdCb,9C<QZ?d79OcKg&EU\-<:&\&P<Ib.&73e4;<)SgXMFEc;
N#PQ)HKOS48>d\+@1G4;+,NYU&F_/XC._];_RDWN8V1]/I0d2AVL_C0)UHdQQ^LU
E001I/[Cb,G]K;[C+dea@We8/]CH3IYH,-;S,SIX],[3Ib[[GD14TNX\,)DD6I,=
Hd[Xdd_@/Ce(IIe,&FI=JGSRMO#,DZ10#5RO-XA9NZ?EQ4e6NVe#0/B;8(TQB[&2
+G:OR^#?__6.W_d?G?LL33&ca_bgGHW)eYJ4>0-@M+J/d99BLf)<KLHQX_<G+9.V
gF,6fD?D^4CBc>_gT[bNC6bTY92K<3&Y>PAf[TadKaG_N#e5PK;YBSg(N?#=a:ZJ
0eeWJ3D(@7&(c?LFI_#f.RMJDF,3a.9&E&3J1OU@gH44eLI8UbHFdJd[;8f>BJER
\D/X\adN7_c-S]bHQ+>B>0?8_0\(X,:1)ecf^eFF2WC0Zd8933<Lg9;9[fE?N3EK
F1@>=MVA:]b6KKSG+4eCYM?#DC]J]->K48FM3-[@?<FE7_95b&(3dZRD<L0Pc1R?
B6U@W(=X>d1@RVf@7:?[\\[@GB?12)Y8LOGD?2>N,_#;c&?0\JKBd.4;b85Gc@]E
IUDHRIXXL1)PA:8.<?G2.2XF&dR_Y?VNRVe^F(55QeWL>#c95;B^A;T,H<8LU7]K
)H;?WBaeZ_WR3PJ>KSdV[.@2dYN=:c;E@G0>+d/PO:/L=b1a/113(?:VK#Ze-W#0
&7NONCEK3)PV+&=[]GAg(P/(O?&/A)f(eXJXJ+0N+;20;C;SQ>B6MQ/ABKD?78Ge
7N^&-<-VSKRUN65c,4fYG/]8=:/(X+7;,W5O.X9ND(=[HFTS@8_FKJN^([>&Y3a2
\1<38W/_OL_1G<8[I>9Z)_FR?GJN<CL&=Q;_\4X>;&])OYKXe#@5G597g9RVY&(R
(7&BgQD_7UZVD.:.5d:YHaR-BA/V[.M;X&^(T7gC5GKN56>HdMD(^LeZ;=FO?TO]
/1a;c4B<ZLS-HI^2JXUXV0(U;FBU=:X#DOAZBN_DA@/^;F2D5XYWVRCN^O^G03E>
:SZ+G[S(3RQHQ5P7K<A^EB_&CdTdVa:1\.@\U;JL;]AX1?+:RRRVCc1&7^gV7,4(
Y/D.&,(&.5YB:4bc)+^035W/00&+f)UTU-V1KLCB1L-+f+RdILa<fMIF8DE#-RY,
NWV#9&[RYTb<e;(@P6?8].Vdg9F[=)b:>@S(?YJC?:Cd2gKCDdA\V@Y@ZD=^eHd_
R4bbVP=7?)bRIDVA+c-W\?bQXNg>HTF;fDb\Cf]3dH]E#)U:T3F]^4KH9)5Z(ebW
=#Fe:^dAYSXbK1MOH5fbW](AY-]0I.)3CG?34@&eX<)+VGC-(1JB8O49..BKM2&.
D8C&cD2_>D9>LDUTE3B]_bHWgM?L?KMT6LOZ&3[==;FdCPV\90Db7;IHV2:O=JM^
A/BYYHg3P5#BK\4OL6PU,,ZECDA4ReEaID.J6=Rb-;Z=:dE>6/Y]YMC5N8<FSE62
;-.C=31S?WB;H^=EGFN)@_3J=c3OLcVV\VWdb,aZ-))&M5SM7g[fW42d_MPN@YT]
O#f&D.CEX^O4L10(K@^?QQE>KU]Da7bF-:V#AG:(9M(F>@3fFd=>-M_1^;Q^2cU#
7RA#P?^G@2,.>#Z,G6fC9DF.#N:HR,B:M>,Y]W3G1XE-RP?:.>,\+T1S/-H2SA7A
K-K30]g27cOL@G0G)D\=#Xa:#,1gVMDb@8TTID]9C;De#VV^RS@OVJ&.F_GPg6:,
#d<9]6C\G2<DHUf8U@Y)P2+N9#KXeMJK.3I]^M<F1^FI\XZ_g>CZ]Y_3De@/L=&_
D5TPY9bOA9;CfT5>G50f96LfaDb1S1?4?[/(^2bI+a&?MBU4c\dFK7YI)[5X1S70
#[8:EW;.F_-VC9dOe\L48AVI0;[:=GW^AP_RO8SIddg/_g^a4FF)NGPXV;G@g9W_
C[E:N.?+M4,cZX/O>QFbKA]XO+5@?AK3R,8\7HUZIcLUVW?60\<<M1^Xa<eDB3QH
7M[O4PGXTa2L.@Y]UV==LRONPN(cJCLZNBB2N?f+I9#WQ(C:RRCG#S\OL-ddSgJb
5\c,>c0(S0eS1fgeFeB/7[QH8T\1&AYH9#08LDeT83+Q=#R?9^W]g9LDLOTW?AaQ
X9Nf?J3_gE\f9=g.IMO6-FS\4#_F0F/\<2GRd]#bWIT&5C;1N=JeY0C&4:gHf(<f
I[4aOW[1gUIXfQ3a.RbZHW2E-(Q==OE9FaXMR(/BTFUbK3N1c^O+d1)RJU[Y24Nf
6H)\UD+,Z=XUK=&<T[:aY8A1Yf]3\Bf=5bO+Z0//+>7S9&QZF2Q-Oe(>9I:H#8/I
9)VTA<9#<0OV5PC,K-OW&_d+:>(_,IeKS/HH(.81ZTS>5CI=1\/KJc6:O?8<AWWC
RQBKe(R(9WRV6Z5e1NMMB7PJbY@+C/?GV7I+_F(c#8CZN8^Y#=3U@)Ya0f:Oa,9a
T5OcRL:9ZDN258:0f5.cY<,8B>QcA:50+)?b+_;1XQ<<)4(BW[/c@-KM-]<QZ/d=
F^J7.?U<-]e3Q#F>OQ(_BA6W?0caR_,3bG2X1Q+Xf;AJ@2C)F\-&4ceUE-4FQ@U6
Zg8)0H?E8^I4R]4Q_GV(cPC9O<6IT;OeOd.?A&3TKLCV-:WF?bQN^_W+;N=/bRB2
O>0Z8G6Xf5ZOBKRLD<J.6></]<JRB(&?@+T+)Cb[bPeKF=&0+9c@+&Z@?9UB13b1
PX2H:H<LS:A7Z._\9TPUGg0_]Dc7]?0.539EA,[2#?2(\I:^G&V1>^<gSGB25SWA
TI>B[P&A2YHf_[D7LB?eK8edEUT(?30Xg6_&O23af2_BKL8#e.M#SYR1E8_,B_:\
I7<aeaCV88)Z04X.,1L>GI_^:A,6;-Hca\/BH74bB90=F4[XX#aKgOg5?L,b-EX#
X0&C#9R5L15-U#X7O4VWca<L5>1gBJ8+2c;GTeSY)Z@.cE/d;7>g;A]V+f/@4BKS
(-,TXQ\VEXB-?UT<eRA04[C_N2T=PO.(6gfQgFaK&eg&L:V.K_#TL#K2[O<)4/J:
4+NDEUe:_)cXE-Z><C>GDPZ#M+/<ZYF./c7&:-Y#aI.\aRD.>SL/WNLT3PE=CES.
.U#P^gg]U7OIM(f68)=e=W;WCX;-BcZD8a(I6OS=&JA_A[1CY<e>_gI)LD3S,8[N
W?UPS<7[=ORB/5LRUG&c\>T(gNYD7MQ2:2V2bSecQQXQ5dc)P1<.Z-2S8C+@UW&/
5;C8d9eOMMf:MaQ?V3JZI99LH]Q,[3R;BcJDc^6LTg.f&Wg=MVU0c>+?I@C_L[1W
59C#b>\,XI9^;8PZL+F(2C6<7SK^RALaW]Gg]e[C51G?6DC./KW?(.6T]dbZMVR?
=?Le>37c##dUZ66RV(>_IF/9HKab,6.,J2A^=N8XG#abfI]ND+P-7M9?CRU2HKP.
<4=FPeV;83C)]4P+B03HEUBMFRaY^0FC&5P8<[.XPaKO]M=^ZT9MQBGO(g?#=D>c
E0(-V,Y9/7VP#(3\A+aS.\4##H/U&A<;dMY07),1RKWc&SJKE>6UMDOX).[WYU88
HXU851RA&)<N0N6P[:<-2eS85-<3(=:(2Hb<acE_.90K1PG/MQB?J<;.6J,/87Z(
-L&^D5BNT/]G:XYdF5=DJFP;@\2W\>VKc.aSf<+,OaE]][17D#97HBOF5f)H-ddU
#=:CN:-LY+U>g/eV.]M?TVL-b\ZDY3S,WabC)=<1^9I29#H=4+3;;PTPQCP_>(>7
<7La>E4HL#R_D7afZ=;1/?2I60eTG@:XKZ)ZV2R6P[0HDKGdW9Q(992A;]JI<:UC
K\EP9F0S:5YV&C(3N1=-+K((PW]6&[Ec/JO<0=8+/C=a#RD37,ga?IUdHa:)XSTF
J<3AJ.<2ZAWe5P^Kd8SOHY[PN15VZK7QV_8T:&0b_:]O<;\CAd;dXX/R3IVGdLbJ
8)P?+]//Z6aEa)AcTKSOD=bb1EKB5SM2Z=8F272A;YC4&&.WVb#C4Q,5\Q1VO=^T
0BM0\@PO[e;g)[QB3FSXBAWa2UJK@.),,N#9I01F#\IBG9B,FU/R\Z@736F]=VI4
QT2663SD2#2)dQ)4UbF48,g7_I=BQJ>#IGEOX2e:2N,F]+<b62>O1VF:PLcY4a+^
H,]2#\1V6/1>I@2?KH-]&;[J+:+:>\:2JIQD;93WHWW25B6.5>^^^YT;RG:Vg?_S
ISd:1@b,3H0,.@gc;EX#7;@e\;-YO7D2b]<Q0OP/#=LQ[:]G0-V[IW4Ab-9JP^Wd
B-LUKELA:,9_Re7;J-WG\\(;^dY5Cff8B@]D]2ID)];ZaLB;;LD.MHP]=RZ6J@OL
0&3A-PbU1<PEG7=9[Hf1^O<U9JE8:D#?);c>9>Xb7CV3@X0L7cWXcdZfNOf5QbW_
EV6T]cCK0MYW)b-,g5[B1DcO#N[D?LC\+^=cOU3[Z/M7V2.[f5#eJ;X(,a65PgE/
FD+QCUVa/7&ea9_;=L9;O]R5AEe5&CGE+06(M?&Q0G87YbS#@c&5g.Bcg-->IG04
+K2<ZMDYg.C>MTSG@AbS(0K+a:(ZPL9]IV&Fa#K/,5DQI?G7CLAIFgMMU6fdZY[1
]X2<+#VYaD>dA(AFJFTb3GcU2E?3EABH]#G\I0bYcg8-eQ^_fDFO5#W),Ec8NOKI
3G\P?KF0K-bSVD^HND&BLY8I^^;7IefZ1?T@T;0g1-^].Sf,6JeFW2)cfBPB6NDC
fa>0\VOHR0]1&]5+U>[?T[5@INM.WdaB0E9Q>C)5c#g,SY_AV;>J=^]P/\_<e-Q&
<TFF:MXC9+7a)H<W9Q(_Od#Z,P>\7YCU7(aE1c(0g)8Z](:14SdT=1VL=:=(:6/?
DIOUbA<Yb(ZP7,#?1VQM6SM_[fON@2<BXID-e<55cdC)7:PA-XPWDRDM=eMJ@T1R
>g@g:6g\LG2CSM/bNa)(ZMCa]HX37b\X.B3V7eN1@R+=+80f1DB^ZZ>cLXLIe\.U
FQBM\@F)(f)aC-A/[_)EUPD.9.8_3=F.,G?65cS,c@G5HXa#I.ES,VMKA7N)D6YR
ISfHU/f9:(5?RU@AIZ4QKT_:DDE)_I,;dF@0M3aG)+=TU9+8;0Cf/EN7@>P9V[aG
VD.?T).OX)_7D:@DJeA=(#Y[TAge&8P]X>b<]_V6+Tf@^ZY<;60JUS#KOe@PNI0G
TfO=WgM5aMa6,?JE(Y#@(Ka^LPT2J[H29(O;CY\;I]7>-:U77+J=8A_4,ET=]:85
V1/3K;beF[L257XYW,_VfB5]7TK\+4N,7c5gJ?TXB?16=3\)CDg?FB]H^K+VDa<b
Cb,CI[9g)B670[1=4P-fKLc:ZS(J^X=g5_aU??QK/YRP_1C8:eDVJ^:ZQ2<8(Y0g
]TB(#LO<]Z5#0L.P..;@8fW:C1.gCGPNc135V(D?BWV>R8G(_V-&a<JP?O0S2>2?
E#BJ4\16J@bdG]Qcbg)DX_(3)XZA1@KE\,EcB=R7LOa:AJ5+FIgPbRW]d6b8KdTC
HPc66TB[Z6]7?DRF^;]MSGY?#+I9HEGcXX[JV#J-]\2;GL8U);<VZAQX9SK+34AU
FdDXA.LY&[SURdbE\^#[M.-<B-bU?D@-_A-K?9Q9T4QFZ,UL\9&RJT^)O?@0e\J8
eYdRC[S-42PDdHA6W##,^G)-2;bf@C:4C>]QV6AL0,D::gb2Cg/WAX=f#@-EK<:3
PG8NDTg1LJ\K>,GIE5N0JXOe5^):K8I=-]G/:7+ZQ7bJ6ddZ44S]#-:/T[88f4GC
[HbIcR#3G373e;g6L#f>gJP2?)a+feM1,.#d54Xc;Db/V?05T3><cSSe7>;+TaDG
LK4;4Fgb(J_S^0A\VHMb@0fXe)@W-@WgNI.P-<[??S(L,.<aN<A9#.b]T[36+I/M
bCY:N_<W0A/7353Y_EdAQ#KSFGIQY^BF?R__=,@PAB.]Z;T10:=gFAK1&<2=J53&
SR.(X1VTJ_aDdSH/O_35IdJKe;QNR;6K^gQE3aQBH)[DQ+9I[=DQ2-#>-P->ZXU\
&a6aVM6AR9J-LU=7HHAd>O9a]+(G_E\7O(T#b=IOF91;&U559B=9D_4),C.W1T^2
R)70@[(<(QTeG7#C#5#b1]I/FT3e,G4FRFN92;-(A4a6-&_gKQ0a^dJ\DYZ=>F7+
_Z>4gZc-8<Wf&]4G;<J^6Cf#H,1F(5=dHfVaKb^S\0f/LL&.JYBLCQ#46_(4HHG?
cRdF09+eVV+R>O]Y#KA0;XL]PXg>4&^gQ.f@Mc;GRT(,;[(+;K/8gK(+Z9^-QVZf
9I5Z8RM79P?84/58X_ZQE8UT.-:0>K3\8B4JAM-./XRC;0ZF\PG_aBbW:]2FQSeH
N[2JLSU0I?d?c)T-L@3S[<b:E6Z#9&9?Pdd@Uf.J2Ea8.SLV1Y\5JN:/CTSKQ2O6
IYH1B@\RRMLd-f\>eG<\.Q9A],CbUC68QNL>cdS?ZCE@RLMR7<,9UW:G0T@cC3+4
0JOTAGNZ?,g#4YEY1--UG:HY<ZON&cQPF\@c+M#IRVZ:2]HVRTYH/].gAIf>A?QA
&#M+WL4We;.7Y\8^?O]&7ZaaY+0:9O0bH:CB#694X12M(K;]&S6Z>_c[;)f]KO7c
I>3KDZa>^Z/>]FP-D/geNNb>:)-933DB;<;^<K_C+62b^W0OCHIMFId_;JUZdaY1
#5@:Q?SO9&/.HXb6W2,<]=[aFg\9G8FGK#-=BX@9#S(D.gEE0@2WgEWQ6V)f\FX]
Q<?F^;f8g4YL.DN]&M@)/GV;6^^8B?+-8:#QW:A<,#QP5/GU,-Ab4Q\X0cE\eRWQ
MT(9fI9g\4RcdL3f.-7>+5f,/:#T>BU+[3(S7,1NK4b^27NdOU?:](TRLNH(b(O<
g)3=8_A>D/I/B,e4^-7Pb388IcLA1MgO6E]OP#M8LY[f?T78P91SKg<P6SN?U<;a
dP5H?Q:<\TG?SD.A9C(K6IU<R/M2Q,5.4RXJ.4#;M/,BG._K-I-+2c=Q=YP\GM,]
.,RTALUWVN4UCM>/S:>YU+VU)S-;SMO=;23YZaWY(f18DT\0-[>;2-16UA,W0MIE
26?:/YME@0<KTO-=BW15YeaRdO=YG>2HIN3::1,<43f=V^43T#eW69#aVRTY/GTC
C5-/XdUE3(K=JT]TW2f2bE?-79Rf>Q9e2RQ\/2;J4Cg@]>OcX/c)03TVQ=&=E+F4
EKaK#E&-cBe9aa(Qf<;C0a?P=(V#/V-EI@M6M5773;BFY+.6Ua46K-+Kbd,4+e9.
fSIgVP+0c-b\E]R^9S3&C1^RRHb?1CGT3W/f@=dRNWO-cE6^\CX:KX::IR6[,R[^
1SA.&HZQa:&>:BBW/(8;Q]Ma7E+.:WcQA4AfOB#E5DBdRTd@R@T#K-<4H6aJGE@2
5A67JGNV51P\Z\NI73675f]2=,Zf+9bP<-=J_PMI=SGYf1J;.RKTQW+^cbEEb&)2
NS2Ae\/;4Z?H2De5KPG\=+\:1=Q^@3=<+3+57GAf8O.E26dHgPg7&?QeW36D]-C2
RE6\996ReO.76_15JC_\2#Q>DH:A0(06L;72GD4+HGU2&.cg8G&^Me23V[gdKfCV
J?]LPW[?8N>6(IATBeVJN0E8[2ZIT/?g\WC6K_de?Te+DfG(=5LcC.QOR_cG6NcJ
7;bEeIOdLEY6PDPX[>,aNKOI2?[-((KIf>)<071EB)K@J4+8BT@g+ZEH^Fag)9QI
&U/(V34S87\#DeK)bfL@1g#D7<;U9@PO7C_OG1:UADBJdQ+G5(B/7b29?;g37E#(
8bDBAH1<G<b:EVVX]/\19We0P;)Za+Q[;;,\<GF(?F:/NgUNXN]/ec[KR+;ODM^W
d[aW8Q:#\TUC36C2RP/&/FCTg<P0H,?GC^LECdHP6(8X^.DPR^Sf0cY/dC6E#0Ug
Gab2U/MG2aU&aC(G8QWG@HH_NO^DWH\]TO,Q+GL)Z>1^WYf1]b9#&c.^TNJSADQE
9OZEZ/DVBHK.IN4Y>,LN1@]M)5/:&(5ZR<<KRR#9DB?X:?W+f?@+;3.fLRPE#7dO
V^?7G+#I(M3e4)]^JdRWPFA//g5?NB+DBQAY^EOP?[1Z-=16R_P_fCS^-dWLG4b<
<)?8>/D+6,6@e;EIE&DVY7S)+cV<NX@(4[?=5N@E-Z30&bT2T.:=U/060+bQfF^S
G\L\B#<9?5)CL:e)5Y.f#<dg994:/a>5]<YG)K(+-O#f4)A6HZ^5=9<9d).EI\&D
,dSKE#.(E:[(4?@3J:FRTgD=.9K18>MY@T7S@L&>/3SC\A<QBU<RJg\I3PdEH&Wa
S#V#E[#,J<F7@_LNZ0MBASf_8:N-[\47c\NU,aaK7/FQ>#3R>;=C-GF_4LRV@.2P
N-+/YJ;79(V=QdL0e2GB:Ve-Y-@HaV7(A;YHQ\eX^OJP-#Dd+M50FC;+^):]9?7T
Y=>)c[S@ccDd_B?_@^DY94B7;dCC&e(^Zd?G)Eg=f<bO?[Gf/RM1ffK&_&<=6QaS
<VJ31Se3A-#CZ@Z.+TeZW>[?11M^R_RM?QF(L6);SS3Ka\J4@K]K6b??5Q,T;bfO
G^YeaVGI+15S_C(_BL\fELHc(C6Y:3Y(SP,/B4YC1QG:/^C[FZfTR3>VUK0b.XO^
)bQ909SIH_I]0^S#6\Ge0eZH/<7\Xb(QP7_QK@fVd@EDYN3Q<E@TeJSF#,A8)0MM
fLA=a0=B<D0T.ePH28;@1Z?[IV3);7ET9^RL=f.@7U-<@Q6&-)TcF0CU<NI,Z^c@
6#L3AD=3Y57/OEU(C?]06QFIZG3S;[@a]fDBN9J)A=;.O/>:]bbLEFHGc71c>H-G
,P=>38UeVeg7BZ@2]c(<G7@6-a)7.f#W<,f_(PD:UbM4WL_#TXa>@(5LHJD_)N<e
9M.E6?-&:W>::0DVb+9>,)+NQ@[:S;@.YAJ7e@7aWY)/;RD9e.Eb&5K9<[8;-#dE
#_c8+8/QNC43GSTacX0U\KM,)A.Z8<D\H[<Z1Af\\-NW-U-AFX26IZP6<3MU\^FP
(QJe_UKgAFD_aMI)FYRCF(&B4R<[.?AY\<:1Zf_Y71:DV/IX(+SIIPNd,7:;&LC\
a118M&DLZc;&F5HbIVKZ(E/f[bc2@&RU@H_KHXLf90LR,#I#YD86[MU8TY,MDID6
=Y7D/=UKRd+E0Y\:0S+_<N4?&O\HSW=O4<C#1Ofe)H.BSHbCf9L>;B?Ncd+6SB7.
a),V7>MEZfZ0C[B].e<H,<(,K_M>b,E(Dg;3R2S@Tf#eP#J0@O[;7aJ+2:(1/R#.
2GJ/2N\QPX179PU6Dg8bAc#bK16&]KYSg<>?_W3\0=NfT-R:5_@_JJI/-0Fa1>PL
?D8J70MXDA;@H.b_J]6AD/1HC<H(@[>&\4eNE0]EcB&87G7[,J.Y^-(989>LdDG>
R_6NNY\9<[@F-gb^dV)JTSK_)9IORPOQcJT[2@N3WR.5Sg?ASK03+8GPBH<ObTIO
e5KAUHV6\=&BRJ]^M,ED(Kd]g<7ALYZ6Pga9C8?fW?PddP7W7Wf[2H5D/I_F\^]:
373#)P)+IA54@@8EN9d9RN]GCI3:B#;AYZ5cXe:9<@:g?AL.RfDDAV[#[OTOI/f0
g14R+;>-Ld_QV8bTQf_R07<^/P@I@BZ-5/TE)Ed@YVCSFeHcdM=;\2M#&I)PX^AG
6^;0\S+9FH:PU7_<Cd&-FF^9aI6[aZb:VI)^=6ZdBSXPa:P1G6ACABc<eGF(734]
[RLRG<9ARK\Qdg5(=P^8GG;&5T^\0a#B.+>7&O#IAP\U;gV)Sb_]Ve90R9C8:HB2
NNF^L2JFE;#LY>IMe+I5P5QU,LP9\47d)ST1B_>^/VIf[K9aPZ1DHcC.3S:e)@;C
LZB>[RIZYaf52(+>IBKFA,>I75ae)693f0ISQNN1Y4^eCO:bL,)I^_/&N7+GaH_P
gZcF1QAF4G/(d/B2cCeRaJ_Qc0EQ5]1FY/V924BK.,FUYXIPURdT@cRNYg0J?ZD<
7O^C]1KY(]57<^2WHTY_+XZ#:)PbO<0_;U7c]A6Ha610fT=b&SULP<ELgW&R]+Dc
,<?(=/QT8<>=E)[W[A8M[0##eLM[\0[^_80be=772:,a\5@WKK.(QV>UZbaf/)&+
+C5-REALKN;ZFR.@7HLOE>7_?YFI^E8.:#[OA<>DN;?;<a\?;/7)2AZ.4Q:\8>XT
(LF@]-W00QK<Y,_8II@ceHNSJG@3b+6:E#.@>J??b)Vc#,W6ARWSOGW.:4,&EZT-
1&3d<bGb\g2V);YVDORa?d-E/G;5geaA>\^20KC+-3M416_KN743b>9LQ_EbRV(>
N&&^D&?a)_>Z/:<OM,4U+#O9bSU+?KcGP:]_=8bPN&3/f6>-?DAb-6SLAQN8gTFI
YbPZ^0[d^H^)eYIQ(<:bO&aJ=#=[R0V+=G@&<4<5G]/(/9&YG(S:Nf#CQLS9eICg
&]Q(/7AXS:.N(6Y^4-5SLKOE\V6()-\;SHZg^+\)ACDY,S-H?CS<X38.5(SA8aB@
Q0KQI>TUDbHSJMU82A6@eT<e/FA=aI16T3C(@<)_,#(C6EG3^Ae/ISY[T4Zce053
\5)&DZ/G5Y+\F&O\\YZPaL/..ISUT^:5#EXGKN_H]>aX\-X+8102YJ>S@@.IJY:4
99CM?IQ)fDK&YXba3+g68F#.Q&be72@U-)#@ag/Q?CLFGT1,[G&^-:2<,<L[GKER
;,ERJ0d05Y59.&aJ.-fJRB0S)=<#LJF4:J]Za3HbBdf[d)\)@FB>&bIG;99gN=\X
bW8dQGDg7GLfe\06WgcY/]3M3U+@Q2O5RNQe.4ICgYP[A@?R+5OA>Q_T&0XJ(+;\
21+#B\+ARF[D.[J1;;1)-8_X@T9BMaWG/GTd70CW.^;f:QCNfDBcbMS7K(8fFU]:
J3d#6>ZQT<2D9,4E[C->Z3_5KMXD?C:\S]5JDIAbK[DA5Z,MOfEPW4-)/40JWcN0
7F[+0P93I?T0eBM:\SY8?Z.IP04.&6.e:DJ<X653UL6)EJ_fa_+K(8>4A++N,Q6U
g&5J9=0+S?aab4I]3Uc3NI4N,K2I;S.:bUJ9X8A&F^?KdE2@(CaN^TPe04E?AZ+=
_7IS;4Bg/B&;b9c?_@]_f[:_SZXX>/:\,DRMO77bEQU1;G?CX>2+WJ^P^;3bMd?S
:gMD@XWBC&I#[a)gL@bOMAC)GeY8Je<M;Y&=0D,CaTFQ116&)QF5dQ?MO/,^:Tb5
A\P5fJA,d#,5MK[T,Pf??gL:VYURVEQd0cKM0Id[1@CY&N]bU9MVH6OL97U2#^R6
[K;HDP7Qa9)gI&@cRfa2+a0CFAd(^G[E+UBF^EHN][R&dP<IQ[[f>Y1D:<9I\QZ)
FYX,WcaO9A#X0?0HH+HUEbUfBP.6>Fg)c0.#ddGf>0#MJ0IAM<)6,eT&be/+PLdf
5&3P#,CC_S+3B&NbZ:=J7,\cf#150=]=OIUfR507)b2GZ(S6<fO\cN6PE]H]8gAQ
RWHT7-L>EOU+I7Q(Y;H/f>+Q;P/I,[FM2ZZ-?@:ON?JVXB?8H3dG(L7.VbBOL,=1
QJ@V-::R1I<ZTIX6[+gNQcWS#YSWSF:bYW/8;:#I>U2\:Ie[bIcNP[:A?R,g2\#<
LS.\,gTPV<ID9LK-8H,U0#WQT\8gV6+Jd#F^3e=Yfa,5>M9dMO<\eSUDXd.P/V/(
H.Ab4YcHDGY5g8<SCbbf]F13H>FgYZNe_:D1\aB0.,PY]R8&,GWc/#DY/gX:GP8G
LX1J3UHH<.A0PKTOAGMOU8gZK\:QZ<RBWIFJ3XO7gANB.]C2H._gIT,aPD3IX-a9
WCI?I^PV88@:O2OUCHg:,6[L+H7(_7;0/gEfUU?6KY1Nd\5AZ4@9NFXfG_eA_SC?
0-?,..DU2P(e[],70f6DO[AR,eO;4P/9^AKBdQO\,Ja,,2(R+c,J(.@a_\#IfB7I
K;?6J<#,^fD,D2]2ccMS(Q4A1IM:FT)8C<g-TQ59&;S^U&3Xb49OV#Md(:@0GWIc
V5ZIg:]CW.6fF_TD(L9IIS4Y7_HH[D2ACR?9(1CP#L/DEUcEg3Ef3+af6L2e.7R/
^\1-Pf:&DO]7L6)\#5H^2.^QAcA?>)B=g44RE554U>PId,OEDf2HHC:eZ8bYeGZ)
VAVHe#Ue&J6;L)JFN\,VQZQ7A3fd(3]U9,))6ZI9F7;XT)0V?g,0K2e5;<Q(EQT,
A/Q0Mb=d<(5f4,Q1-]Nb[MRM/&WR@-R4eA08IQ_\_eDf8ZEFg=b?:<VW6OCT)6Y(
8:_OCCbI,JcIEKL\@6c#OT,AOSEIP>VN15c:,:BbVG4YHV@Ic.8I.N-.W/\I\T#X
9TFG6^J>^5e+=(g2QTQ(BdWRIcBVI1F-8,D0-]/32\+gg1FaBZL\[MSPBb_9.AdP
e0?Rbe1+=:Z:?SWY(:GCBELX&eBaf)9:RY59J&(U,(&3XY)8ELTF?(R>K#EJ]OaJ
WDRV]:d98SXH2LCS#3N7&ZJQb=\7YW,PKAZJ73bag.;PAM5@=5C\B-PYU</P0T\a
;?@YII_5F35@:W^98\YaXSRZA&ZQ88\V^FU1\C6]PT8Gg-Ybf\W6I\Dg6QQJNW#M
X,[U&>)M=#4PFTXED#d6[B&e::8T/NaTJfgXG=3N(g7\-GSIQ,JKIRE\Q^+GF]T5
>-Ue)gaZE\8fTKB;&RIYVeNS6;R?&M7;6e=F8OSX#/8:,J>Rc2+(WCCR-f7YRe_f
YX1KbX@fJO?)f<bMFHa+FFJ#-aW>WH)Ta#1L@X=#[(8>d[QCe7),Ifa3HO3W7(D[
K>aS-##H4Cd4:E@J<0I^;]F_XT]-W1QdW:1E1H,#<I5(H=;H5(3W9M8J7F>eAWf[
OJ8e1d^g]g:6ZQA2M6f=1\e=3N0(d#:d&?MZ?E<QC\fNN1C?.)[RRKQg3;I_d/2Y
UgXEeW#Z;TgR0O7]B1_)99Gb[8<2b&?eS.MFI04]8+E(;;9ZHO7OcK4<^O;9WKGM
KWgR<((g_2cB4d.3NAPPg.cQ=]E3J?0?Z^AfK(IXPL.BFUPWdg]#36B1,VJ[c+Z;
,=P2?Q/]-BILLA8RDU6g:HcJE-1BD5AM86GQ.4]2HJODJ_.??5@?dZ+P@V6UZ+/G
Y<MdFV=9f74TYDY8SePF;M8G2N>O;U7SPL2@]aF=Z&WaN2ITMFAU>ZLJ;g(4U.9:
&6AWXG2a=EYDDARb]V[HF=c/3=-Qd?=C/5(d:JO9];)3#OLW_;KO7G[I/,(Lf=.I
B06bg@[:(/g@CN8ab[H@#KC4N=Q.g1ZKH[L6;^dIc&@^RSQC3e8TYM<B9#DDF(1M
-B-MU^I5?D[(BH\XZ&3>a+FC_EfAZ]ee]Q0;:+)OYXf92@SU5S655[3R-?PFcPNN
e+a8R7NJB44_2FTZc/VfK+(+VeV-0E:\aDWd#83B>@B6/]/RC(Se-Ff8&MBY#T\7
bJb)HHJVW)<8C(-2/HFI@PPZR4?Z>YNT\QCZZb^eO_d;3-3f&9ZX_B+,6bEJQaS<
65?Of7c+IA^;]2SLZ^9d]-6c+Qb(,M<A?d:D/5Z89:Ee-,R[bC+86@W^2DRZHRb(
K/;bESQ2f&S[)18@5c#/JR#,-];#Fe9gKINT1-I2/5PCY/>,L0V_,N>;H0Pc&>\A
+gCNVZ071.CT?AL^TCX-QG,RG1Sgf@8g?8_SR]dN^</RU>+4CA]ZBD7bVEK^Z,GC
N+Rc/4f]VGIB0N\f(6PY@=[GYM<d+>KAL\@-NT\SF47.5PU&A)M78ZL>V9=ES_;&
:@649#@L[2)5HN+cO>fKO<_]AXMd07DGVC&JKO@1R]4_-;BKc-M4bL=TYR?Y>.8Y
C8UZE]5(-.[5PB+&I(,).S6/;?)Qe-;D4:L645#(5<N(U1):6S4L:<[0caP[)KG?
<Rd^[Y0ccUPEAd<G2_F(M(Bd]Z)bX@\5PK[[IXE,gCa@/06V+T3YbC>V,K8@Z1Nd
<;D,d7F).=<Oe6ZbB2W,L0)N,E+JSIPUM:B^?7\Y.L>ZZ^VIT/#<83N9Z1^SO8#J
(WVC8BW\6-OSfBdO9:FS^AW3M>IA:_(MAS)K]SA1J.LS1GVMa[(B^QBC;)WF9=Ab
0^3\SE=;<UcMcBWGRZW>PRCdCMg1VL:]>9GI?9A>F@(G4]B((>U?0-Rf4XXT4?Y\
<,3]1B,[c@5ee^DaUPf/:HX/[5BE<YDSC80,GcUG&ReD7TON2;aMUU/)4H.\-Meb
AbdH@W]d@SE[4VB31]dFbd4#<K\(Y<2)TD+IINg_7X<;62]CH,Lf?O/D:]TQ\DBO
>GIZ3.IBVJQ>.e#2.PeN8DM&QdG<.&J4]a1H.N(9:U12(H]S)c@:IfM3E<&QYH9T
+?(d->9K7Z61N>V07.eL_W@+[dggGK<7\e[BO1U<C/c:CTN[7\/-^3,Y_IATObD8
dMGAL1<[_Tb\@EEXdOKG0C];N#;&KW+d??<ebF960JK4c)#D[afS2/+4YbHg1SRO
;@[;&\2KS(0]^+AIHD=6>>J@cO0D.XeOcHWWAT4#,cIX>RJK+?UMSD<V>32^CSJV
fLH.B5]X>?N2eIR^SU@@K_EC9QH7/MG-ROI:ZAU:VH3;a=@c5Lg&S8X@L+6?&R5X
JU#-_/(Odf=UVB4^DPBEP]9/=aB7bZGPK#TN72CP#WXF+gL<Y4D1PF;^@bH^W=^e
\#.2a&3\4[Q](KJ/a,5:833]=UI,:<I+185_RHX+ZC4T2&F3[.NAOE=B)d:T()#]
BFVHe0Xb4-L#HU@_fcgQ]fKa)W._19:.&6GXgRV(4P^,HWH;[+.]#NSHC+#Z+e6Z
6P=U#(5@IYe6Y^SI_>Q0.X#+WV3RK/&A;?0D/AM#^YE,_R_b=O.A)C:WPVB0QLMS
^Q2->OZ_:@:[Gg0JXKVJ98U.PG-CM560]KSgAF&PF&EY.CB:,XE[S9W[9[?F,=0O
T_FJU]<gd<bP/Gg^>d7Ic:WL0<&1@YT;Y7/(c^O=R7e)YJ)0RUg_OH(M8d5GA4I&
1cD[6NIVIC?OB,4P<#6K6(-)=TbfVZ?U/&J?]:/9\>MKYgT&?#6^]X(\_GXb(CE0
D1b]4+6-HJdR]@e6._G3VXR:9VREU#/\REP&PAP,gS2f[OA_[<:Ae?]BMC>4#F#1
OJb,^CL(F[W_7#.9&b,MN:/I=Ydg&0#?,W9e)dRB;fW4TeL.CBAD[VUJ.:EJD_5O
Z;7XAP6_4_3Z:B80A7YUaLKC]89?P/^=>cVa.eT?]g#U;b7J;@S1PY)784c<(^#6
JYG:dS2C^G<P(;Kc^;=((@OMA^#Sd/@T[FVS9?a872+?_9,)-fF(ORb1GD;b<]F6
^,8J-3=CM.<AIIc18J)fU26^[:=Y+c.3L3S_HK9\3WcT/0X<OFb/YUSdg&g0E;O2
[+0aK<K>7c@?4d+>F53Sag0\H9WA7E-FCA2OF_8/b[7/a=88X:.FVCG4^W47A;23
T^?3_14F.AXS&SF)>3\KRS0+K=54#XNA2_=aZg_GEMQ/7Q8;H?M>=_</.W]KTa/,
/:Y7HH\742UH[#-_-^J\#(,UUZ9XHYHZ;GSFD;F>MO[2OIVW1JXC.g&>O\T_#@(@
C@+=W/&ag/6EW=2Ud>g9JD\9N;EX^QJ0BI0.D\Ja#4^_#>gPcG;CREQ3FZ?LWgd1
0_I:A(-HeJPJ/F4Wc..P[--?3#W>&_YPc&00a,W<8]RYZJC-f6U(Q.a)OLGDSZHX
4J3]g8FAcI]Z+NZG-=N6;Y\f,_?eX<+A<WSC[+J3+9f-Qa/:G(>+B+,G9C)2>?N8
RbGM.AQ.^?\Pf@DK):G,NP[b?8(Y.K-Z)K?,;?cG9973C9T]32XGK#PV^>VOVGNE
+(@.T_-f9+N&ebH)-:Sc>2aeQS]L48V/A,CL;=TU1Vg;Dgd6YBU\>5=1V]d[H0J1
Z+,EG]2TNFC3,&H86VR=aKA0fE^@V]VPA6P_4_MaaYASRLRT\,WgIWM2?Rf&YV3I
7HbQ&8-V0f#]b,@Ie/@/cNY:MZ=&7SfUB<Q9K+#OENAG6>]S-4+QFR9(-P1FDP8d
DZ2/;Fd)YNJ\:48W^^C@?B+g,D,6T0fQ?:,CNB0AVT@;:&T>M1O3>Jc7;5#2b/P^
1@VG)758GJa[6SM4>@b/2g;Q=YO7Z7O>RNUf9Y^Hc>[#XLC8SeQdKb[.-64A7Y)4
;BgA.6O6(M#?:)4KV07A/I0[\1gfb&(8Xg0D1Iaf3LC:M_Vebcd0IPJ_<^^=RPNV
.W/S(C2GNad<HD.(:/@^)K58IgONW6S[<_])8>Q86I.aEK8YdW;gM[6>TBF(EXc]
<NZfQ^D?@56Z[YOeFQ6dfgg.3)(2LN8d,N9DF(GIXJc#^S<1.?BPg0JcR;/gS&;K
aDXP,LKJPY5CQQ)6d<A1C),6W7YSg>SM3\-UXSPG\)@<#aTL:F<3=VI]F8&I@O]L
PV5B)L68F>N.Y_Y:&cQ/XJ_5W^bGdT[8b-P-cFBO>4,^1ceA8?7PIIbY#IIP5L0;
bbMN8?J2IW^PMKERCc9T_e1T<NBQW(I@9IWIJE\J32KRe(9>#<AH^2BI-A&&caB@
M3_9CSJ\J8UM[)788Ha-&8J[Q11@+27+--#HX:dD2FZ;<@G0[\dgI-TZGPP0=<bf
7I=69IVY3T??8Q=(YRKNG=,<W]1-,FZB_UIW9#,5<VBX^9YL5#<.XIMZE_(Oe30a
5CM>bIXeQTXL2A5I)RX]BFMJLPZ49YC82b0?S//I&D^Yg=0F82/K=,?d7,^Z4+9(
1I:IeJL2B38)SF:WF)ae>.\.QT-WB.8gV;EJF3aN.;?B7B#g=#D<^0V=\?B[.)4c
IIS/BHZ;=0]&dD;[-e>-A9a[TC5J_9UaULHM=RDH8K[e>d&\,HeL[OSG-5D;8H+T
Q6c8g1g\,&-.Z,2(U\b.e+>C0,5T/cU@-GfASc0,:GTR^C3cd+dWZLeP:eXg1NB=
(Ea.S3^3c6Q2QZEKL3+/N@T=BcMVO8ST<56Bc+]D3^6IgA[.fg)PCB1,\H&eF,YC
:)Lg2NS3]&B.E?0:NV4a6cXBK<1Pd8]8[;6,CY-,AKa5:O4[f1^1@0[/I@)2PG(R
E_,f^-W5RE^E+Md=+N[V;5Vb1W&9(YA^8AF6\J.g4C7?N2bOD:/G:E5)VY,<d:b[
_2_0^b&-7<Y,7&43&<^^H?OJ?^6+8.KES2DWF2P#O1Bd7:A>M3JQF-PHR6LAb4^Y
:fVG#7Q;=LW=YV)F+HK^7XM;aH\f.<8@^YAI:S;#MPb;#S.0&WCLc;8.<VV=_,4L
dW@C6(:U=2CN+?YHQ1WC.A]bF0;^2;]\H(M]a[3Qa2).gB:\Q63Tb/abZ#F+NQ]/
]OK^J16/CH]2c\FH#6G\a)?DY^]98P4F[2A/;?@::ZJ(e6&>B&eW;Be:QdQ.ENWA
;P69aJ_U^W#W,,@TVT8LB-(g7MT3dGM?6[:PPYIW:\H\(Lg\8Zg?d;@WHbJJ7]4g
5,;OO^<d]N</)=X@Z:XCS5A+AV.RC:D9d&Wg\YT]S(:-BSA.&&I]VHf\(GQ\Ufb4
)@H5c-EUaYDQOa572,ML=G?@BL+bJcOH]8F:dT-JEYCRWR67c(C1Tg;7)9&VgE^e
H^Y<bTNA>)Be65R@W:=NAXDZM3Q\^I<QTI<V8&ZK>E.>PYITHaX+67?#J;J?U7bX
5MbQZ]7#b@>bFcb)3N<N<DCZFN.XIC7_WJSG;T):(\d0H^GH5g:69]FHY4eC1RS\
6TaQe&QfG]R&AXGFH0(U/F1J1Y8C0BVe@]+O^P7Z-N+VCF@A/AFd3[MR_6=fQ)F6
,T)YZ)ZE;EA6ARdGPKc+B\g\V^J/XVD#8aeN+.=Xg3:6_-5R@;QV1,2<739B17+g
ZXUTeO^8:KEH71_<MfRX#&XKPf-.e7^KQGJ4dJ<1V_BS(If6J3-e=6bf32PCAe[A
6OS-+gW9Bg>ZWRaKCG6O0-ES@aVY<XOX/Z5<=cULPc\6b7(N.JR;<P(8,?W=4:F9
e]fC<gWD8Ze46I9+SH<057DgbZI.RMFLQ&Q1:VB]OX.XGd5)FVT3Z0-K&<c5:3S>
eCF^<HP_2gRJ^&WTg(0aE7:S-7534,:Y?:c;6@:Ra<BK.?UMf;Z?@U4SZaB6d,fc
ZGF[K_0_fLZ\5Z9XY]fLa2?KF@+^34;I]D,](AQ)UINX(,1#1A]V&#?JBb28+A[J
>21C=^a6.EX\@]56N<4U01<O7&(VS_@A=VWTGfY@g[SU5POY=^+^5#?T&.0]9PP/
.2=b&LWP=6+SgVSOXYT:Af5;]IL+P2GI?152?a^YHG&/(_BU3[J@TI\LYB\:C+P#
#:Y^((1Hc7EWBFM_M,C;AJ(b;M]IWM.W[&6KLUZ?MgARMJc,+E7gNV\LM=fc69\6
7^)]VCE65WOX-Gdb(Pd&LFR;CM56DegHeKDFRQ@T4Rf;Y)(XU<J45ZXE<6f?^PFG
1a_e>baV<B8NGON@TQ=/1_:XA]C2EGM)4XQ[Q7c[#]DP,J^14I]@ZDWA]LbLg_S]
RfcCXKPQ)Bc>HB1&+#COf>\D]&6Xb/[Eg^(6&_Q6TUFJ=Zc>&/:JD.^JXKOH)5T;
NAA[]OJ65XG?&b7bO)EH\Q/KJ8)]5]=>R-GD&CYT=@IGb:)P=8-a)(__\V@[37(J
X&5P>5C?X]GOTJR;R=cIZaSMMd0/],>]J_P[<LN.\:S2g&8>GO\,1C[O[:>LI>P5
eYGN/+#)_?2YL<(?C=JO2e@[=U<N\dZXdA3)EW#<9c-.4VJW\RI-_11)#IGcbJ&-
4(Z9\ObAOIKKVb>#F/4]0O6V>?Ua8=CRR6/4E3E,+20B_PBEf5(S4#gK-L8f>EL5
,JgM&W63;+/Q4BfA56b]b-gGXb83A]V^5C.<=7(OR[b>K;[#<[2C8SG:W\/dMVaK
Y^7S/ff)EW+gP^BcB1-=V^RKNS61V3a/PX^7,;4MdXcfG)W39L(<W#@U7CN2V98V
;B=Kg.38d#:ba>bZLWZ@#B9(?JdBK<eS+9),,PR(]3<Q_Q+FeGWcORUWJ&egZ.K0
?Hd,ETK[d.US\.(_OE,H52@+H5O&9V;A1H47D)IJ,(;W#.I5C5+;^9(_>ZG2U94g
4&IHa(X5<L,7[e8Z/IANCfaF+QUK=4cJ81T>3c.Ld&-;JaeMeXQ;3R>89/.Ue7Nb
OKBgP0OBG09P\0Y^=-Z3T;OBAbT?C3FL/\<.]D.dac<U)T/F:Y>+F46=/Tb]=cKg
+<I^\<4AUf0&VY.6&gB&MJCY[@./G3aYWgJU[+3VMA]S>1d@?80^Z3[O?IMC;OH7
d6edZBSEZ5>I6U#\UWCHNM2B#P3L=M0/)a<+0&--S,HQ(#cU\RAV&AR\b2Q)N=EP
_UE,)R-g(M2cC@S71NBc]?X5NUcPG9cgPY&>&>b;@9_33?=0XEScSS[+GfC)LU\e
[Jc6Ff0R1gB06@B@5,f4XE@]=8H/^/b]=@;G?JH;&]7N&ZU5G,).ATgCG8[&&;^e
bFHCGdO][U6C6)33&+WYIa^V@Y-VLI,D(TaI4Bg6>#Jc<3SUFN:/<gTZf\B?3+X(
+eZ4WWX<_PRO.KZ)(]]E::?K(RY>CMR7BA+?O6XRH[dgR^SfCEd@U#&S/^@7GD1C
Cb0W;EY0VPc/7-C21@;4[P[8&6S(P;F_J^S19LH8Pb33g\7CS=ZT/AZdM\PVUSY.
?P9>QQ?\(R@GWZ:7[.Lc^VICSRO#d_T+<_Zb0Z7FaURf&HL-DJC9R5MO&IZ=6CST
US:c)RPUAd],Of6VGKfQHA;e]]5A#5fF:f[0aE,D_N]:&<.VSb97L1.bGddR]4_#
c]?O57X0.ZM&:>G[KK/<(:/_&E:BF>#K?[S=>IE7fY[/K2&2I/UA>>f:O3>cS@W[
DC(g3EN>JIM;/<=\Pacc92AD-gbaN(f<2f&#A<eTSXZ\3S3>5A@ZGS:BMgEa)VJA
NP;BJX.38PN(?&>>Kf0-G24F)4e/W./We[6?-FKM;0NE;]VI:8A,DVFOfL[cSU/V
)[Sf38IN2aRW=/117caL(O]/OAfc/-gJ8N333/R9KIM>Y0c+bY1g7Z(024W@<HZ0
LUR;6XMaKI.Sg97=bKaL(K1aDF1/[9,VF3==I#MaY\A=_LLSS&2G&Na9IabV-+>a
.8AX.@Kc6[ZD0^Kc\L=F3KcYbfT\3dM5McF=,Ic5;^(6OVWW6IgOH,D\3R>A>(/M
4X;((9D0bM4ZQAVHG\,MT+O58HRWYe[5)YP,G7\4KU5&5:4Ke,CM67-Y&e6.A<.2
;,II8CHY2cF:6TR\LQHG<Y.c=2@TR9J-@+Q(-S]0..F&@C-7SAP-:(f^W.b-E^9R
Z.ZPT^\b?#Se=&a:5;P:REfJcQ8f+d-C8OTN^bUC@Y)R7[O0X]B&06JL5:_J]8=2
.C.\#,\5_P+A3)cFCV@VXS^2GV=6V?<\N(.RG+1/T[,AH=?0F#YZDW@#:5gH9.<0
LTQG6CQ,/adN61,V+&+g0/^:63^COS,:UaLeA]VGK(6/H+ILUBdg4U&4DW05VZU3
;(dWK>f]WWV]&T=FWJd2[.N?1)U[,R5W01-\[,=G_5-_@bPWcRBBJf8H?2gScTd9
7gDC:,6_Jgd/)XVND6SH58.V/gH@ZMeDX<;NBDN_B/CB86X#X@4geVC@)^PX8;TJ
6(]N+c;5]8VO=T]^##[Y(OQ@e>[_/7YWF^O/C)b-eDXJ?UUdH6_-WTUB4fT]a\V#
=;_M80b(Kc?Vf/^D++.4K93#fX0[(.]=GEcU-b34(;aMK-VW>)P_C+ffV>V[[Da#
G:I@aJWD6W-67B4&8?4)R[9>]5Yg(;4<5gfOb0EN3cEGMbQ9/U<7/f5f8D9Q:-6f
ef\D7U0>K)L&=H:dc&d0f+f]a<9383a=H?:]Wg,gN#.Ka2,.7]C[gR5(-I+3ePO@
cU=ad><(^^U-Q0JOKc+gQ-OBH-,;&TR^B-G.d486d[T56JJ(+Z;-LQB)ILf+TgHP
HC(V//Y_02)>BX?TAS?a+_We(N36Y>E=Ee1ROL4,5C=-d1C[e.PJS\F?)EH56:T3
3FHDa/\9eV?:P>]fAgTA0Ff3J6gB8dbER.HR=A)F#3f&MJ=NJFAF:9>b3MULW#^K
PF#e;V/TU98<bggR,Qf4)W85@-,_F>a>A]Q:1W:C9TOJO=/L:];^NU(:(K8&^0TU
V1F8M0I<a-d1ELac:)<LG;ZZRa^L(@VS#CfaM(gK3J)#V\1V,<?/)dV)YOEf.I-@
72^45JGXNY<#SU0b)X7R-:A1.;EY0Y0Q20T:>D_f8?S/#8EZD9gc]aZaKF[GgW_[
#Dg(<J?;-[>OeegD?<4U.@]H@#XNN&6=1;J\?0Z@UY7+G3AI,JHK+55YC6c/VT\V
QN1MEgeYc[Ae2:8]b<eWWJR;;RF4bQ3\&+6;QN(9#OF4KWV^S@_[;G(DR8Zf9=c8
^YI8KT\#=VW>RNZ8-W=J35S[TS5R0+JEe1BJ+BWd\8V5TOQ<_1Ha6?2?=f;0S2Se
74KMV.8X5G#a(R]eBZ>WLK5]+FDU78QZg(]:?4e?56(B3?D7D4YYLI73&D;eXQ(E
@O(HI#TA?[Xf3:g?A68&+\G&7?9H?,cIb:OGF.BGY?\T9&U>K_X94=e?8)Qd@)WT
)Z-#6D2bBCHLB_P?KHF+KT@bWC.Wf1<>EG76_cJIYGCUP&T=CNBB4L-###F?U,6\
Y3LEU(6C(3GHg]ORKAdCR[HPZ\3XaG9ee)PK+?]#G?+?[BSbZ56DUYg?a,@FH7I=
I56?US-Sg&9_+F=6)1OfLKWYcJO-M?eD?@bF:-.:UG_OLHDEHd+=UL&#K9LNGbR;
R]55X9QdTJF(X5DBIAJE-74acf_Q_8eWC8dQ+N4G.?SC+M-3dY]XgF<-@aceZ:=-
B36=2\Q2H:f:O(Ua\H8,3-CfFDXZVH>)CFY(UA1=XZ9Nc_a),HbB2@:FbC^T1K>_
APFbRTTO+-c\FD7A,]9&B_0,QZ.C,_aE)QP-^g^VJ+S7MJE/1V;@@8g@1EWAG7Zd
4aE0?9/J,e0ELQ#eF_FcLFJ@&=d26B<L,_)0C443D^^?5Y3H/XO#8N,dK8X.T/JE
<+-6XLb(09K=LbW.H;E\Z/R>=3X.KA3IG\#KG82<<e)=,@+ND],b/R81SH9FG+6T
@)[c&#KH6Za,g:Y@,NGC>NQdP7-9LN.@U>FZ5,,4<e-TUVf6[1(FGS]NI,&cPW[N
12DO(>O;F;7SY;b-P;3_65V(c(TZTLObOG1U^QKB:)e0\#+.WVKe,#I(K@=S7Dd(
B\a_]]ZCd;d/M;08XfE_+IDA0]RPRTK5:6R\33,K&2Hc7F/G^><9UB3@7.fWHJD?
4?E\;Q-)WF([P.?270Mc)H:F[QUI8[;adeDfW&b]GYZAIM82,=d1-e((#Z6W1OS@
\f,SDR0/4W6F/6_bfTUYLB2gXJ12Fc-[#6B=DP9YZgdbbRR9F[A1>5FD0W^=T@97
e=D3Vd9(eAI:^5<<_=54M]aYJ3.Y44ISWX41.#S26cb-4CcKD32XU<c&KJ#\5JXR
MS>ZT<^^+O[d,I0.c<:6H@fWVU@.7=6>Ybf:K>_9a2B:L(cC06;eZ.>aR.#b<](]
GX(>7FNS8T+MeWb/&V>f(Yc@YH5AFe43>Z#TaD=L0?YO0>B\a+#BM[7/g(93V?1+
4.LCR.EL)+U^^d,XB2^8W@4SF(&NUgD=H&H7:T5/@_Y6.9K([@d.K?GA<3J3b@K8
O0g-0A6E#;1\HQF7MTJXdG.2-;RbLFaJ-N@B6Lg^45L6;E<9(=K9_TJ<(P\W/c2?
g^XUQB?+WCHUX>]aJfc>=f]]A9e4)b/HTIP^44QE;IZ.8I.R3/\YB5KVCVagIdS.
L/N-P=]Q)IJXb[4DO?aFS=><AR]R>96A=ENBQ+DA+1dFfFH#YEc^1.)9/&_PR<PA
A6a<)Z(YE/:_c6[&BAY^&2D(NTQ4TJ,U?eOK?S;(6Zb859e=)E/W_#>A:M)[R(5>
(UY6Q9g@RU1HSV^,#G5,)>0cTBU,<L=F6#=J#X,/@<aeYPcb8LE?gX>-GdVB2FV#
5?6EP^^FgHA:]T6Z.Cf1-DU#Y>=c0B],#7fPR9aK4D\P6@3-,Z1I<VR7[Y]aIXKb
.2?:[ceF7E#4^<5>U>dabJ7[e0g?0Sf^b5+#dX,K1,+Z_)969959:MR,gGEZ?=#K
[Q-WH/-BAbHCGU3^aC(WAJK\T37,3.aO.=Y9[[>E?ff43C[C-7#A1(L.;bX:Y58V
#a\#:PMgF_;.TM=a:e;Kd/\<J^O8AD_Z\^@W,De4UUXAC8#CYQgG_</BCY9EOSYE
a65SY><?O@0-Z4C.M3_8WOYB<#+?_dgb4X7@LGbY\Y2e[3FA+@Q]aaE^X5/;Ec<_
2PBe3V\X:VLCAff-1P+fIB5BB.>J52a^AWFEgc[,RM]/\bS=L060B.547Q7+9(+V
ggAZE#C[CcDCUg_GX?Bcd\:TDAT;.PO6Lb73R\+A(BNR6ADfGE<N,--U_]&UHBO\
3I[Y4O?(aK-G7YY.[#E:C][7^O]_d54Gd+2a[);_ONZc4;ZR@:O.ca;(L;Zb(\M2
_AMa=5ET@#]<-8eLQQXfLfZ&DMcL2EEOD220dY=?LVOc4N9f(OQdd@@(AWW=O&63
b,)2b^,A@#72R<^-H7>;&\Z&:f?T#L[&7a<I_&Q@2TVR=dX(IG_1>4\ee>;1g7L=
;[\WeFbc=KI6R9da-QC#-:@F7UCNg]IYcV(TV5a:a32<KAf-87U=4#.SNc806P-U
<<9;@ZfP3D8-X2_aLH?_cXKF:AaB(WGg+_Ef>eBIYLQaDUB2P1[2=1ZDFQPgS0^;
MGYZFUPKJDH@(B(5SA1Q5LNfO6;5Jc/HQ4\US8GZa6[C\abZO8DTFI,:_aLB@.4L
DF;-<]]-&/SE<1B034fNQ2BH+O^dONY:/d_=\aD^UTH,.#]>DI[cP[c/d24<UV+A
)?S9C1PL7)V&&92WWY_-^Y=\G_=3f0ZP+M6[B<6+<gT4e-?9PX7fSQ3aQB.;3-^5
5]/AZUW[E\8a-EZ=;9L.TNeDO_#SFL9/#JVLGXSK-VP[3[eDTV+D(#F1BQ/FCe(E
S,-b4a;HCJX=U@.bMP@R)/0P0Oa)SXg)BQdTJ5P=FO3dDK2Q&;BC:g.Sg/[VFQE_
KPG;X8WDL6QdZ4bEHUVON[-Mf?aN&N_:DJ+RNCQEaW.Pf1L_Z+4Uc<9OP8;.<S;0
?ScLL=0d,Q2O5f-?_\OLe7@L1.aFB>NGAT.dD>Q4.<\38Q1[Q08=5:]\N:H8G/5Z
D&N32,(U4#Y>_5J\7X#QKY6VPS6U:Ug3.Ib1eH[VaJ-VU8;,^F#V.,:[g1)J3O#@
7cAN(>G?g476Ee@fFf:2M1VdN#]T1d99OZI=N>7BBc36N#VZ;VWR@G)\FeSYH@1?
Y_dfJ:6H+X4_Y3gHRDOggM]<[,,68DLQ6OZVN7UEUX8/)R7KdF[a_S)3;V/O1HAb
fWFO;@#<7/1eS^CRK9?767?eA=Q.1_R[LV#77G@I+bS++6f5:8e?#=Ze>D5MKK+D
F[7e5H:b=(,KQDO3/\f7J5SQc\&7a0TIe(cWW\#YT6P2a&Y-[P,PK\IT:LL=4Efg
f1^Ud[+J-^5FMf;N\X0A29bKA8IZ/]g@d[)Z&[bU&6Z3&Y4<aFKE90a#fR(?X7Af
.?eDL7=77=+IC)AV;eNP2#)SYQPA)eT-7FTG7#[?M1=9C&KP77Zc@&+&SN4+eU)Q
-I,QZcg6S#.Oe2K#??P=RSUI.,O1T(E_E+YVSH&1)Z70Va>9\gGJXKeDA+Sa;1d/
@aVeQNXKIP(R_UKDdXB3-&^-G+G4T953:Y-2/14:E(X32SbI.CLgW?_,^KZ(5=b#
\:-V(G[66;N-dag<Y9gccMB(7gB@A0SH_GSf4[<U\<R)c40d;.G&@1M^;^1_)1;U
T0:[cOHF)=?^]FU?KOP.3Q-T[FcJ-)TN1L;@R)J2B<Waa@NQB_:W\MR\R7DZISLA
>JZ,b?:)2Z?a)X1(YN5Pd1:1&]XW1McBU:D(>).;JY2aK(OK[0FYMPFG_8T-A/YV
8N@(UTcML0+-\MV,UI0PKQ^U(3-XafBF>SFU@^,W.gfHg8EX&g+1:J[C<)>>Aa&6
;&3C8GW3N5-,?J\.Ig^I:d&]MRJB/73OH+]9I\T:FRFZ<@<a];RQP#2K\a@fXGHR
L)=09Q\FVbd/SPL3F=_LeKPD@BJH&SX61DK0Q4L4f0V#CPK/6643g;M38>8ETBL2
f[3D>\9DO<HD^?=;HVDETRbG_1_g;HKc_M9Q=[9=79fI+K>#&.f]-1&@?L1\HdR.
7V\2.XOSC\[I10#bX4e.LKAL^?E6GKKH(AcZP9X,Pg@e=3L+^d#OH(E<CLC)GS(Q
4./?(\(E5[Ib8+&[XW^I8H]\a0H_H89=N/LZUG5HZYM=N>[WI2-0e_85\:a@+Z-1
.LG4W_>fC+8=#S1]ILD3aY:ZYY52+4RG+=,Y<\A#^_[@4/NWJ;GNK=)M3NS]3g?=
g/H.\NO1\2.7Oc0C=HBg/()O.(e-8Fd.H9AMb:gc2DfE;dJ:_/DA9/1-28JRM-A_
X6.O_[XJS\Z3eEQd.[(aaBRDK>=Yccgb[YD1@;T7_&-][A(d7#7KXVX;PP_)]fC^
6<AWf79Z7W++;FRFLc7WBO]VfcBK68=#0OC>gZEA2U9b]036\H<T,ZU\8JZ4#AgI
F0(GK@)M(\)KDNcI7^VQ\V53G0\58W[M[D:KPVI3-OC/64.dL]f,+<PJ.3N).SGP
DP=b/P>L>Q_fGH>.<O[)Hb5]>LQ9g_W#02e8;WKD]_X;5&-aaNHbE37Z(-PVML77
^BX,8CCKIC=]eJ[,#NNBA;,Q)SDC([FSF0Tf2]Y6:NR&[\,9T/N7/&Vgf.S\?ZA,
>d;-bD\O(T#0d8=aF\Fe48AJf57Zg+@08>#[f=QF]6GZbHb-Pd1H3.L.09RU++>_
fO5;\8]-@3?EW(8UYLZ4gO>@:1fZ[/g&f#^6+O9,2Mg3c#X(#42I2I1AK/9\Kb\(
I;H)]Zg(=GHD_J8LggN^JF>QOea2^3I:#&7\N,V)G.52DGM.K2Z7F1Ag\SLb:<>c
&(P4e.f[Z5G@IM=CFd-]G04Gg8@.?8ZG)8N6[?>W4-]QTM9B+:QT2.aK(eB[QQ@B
K+[?TdF,NKY_WHCU1=9W2ZIbTe8]b#[ea:<YY2e2+<?:fCb5^6:Y9-W(=ZA18(T^
b2C7PJU6?0:^7d&;4F62#M0+PATZ[#1G>b1&.U25^<IK6V)G,O;X4P;V5@LZ7K\g
0BUE/H9<bQO3B<LX-II9.14/<M\3<XcQT2e3F@;#0P;/d_I=6LOgZ]\=,Z]<B7cW
-7H83>Y\)C,5f&aIG_K#L6c]gG7P68>TI;;&g[+]fU3^UGbEe322.c3LSC;6X<-E
CC8^T]+GBV(]6U#W2V7-Ge=8Lg2_]_6B7&bd](.T(OM-<dW\)Z9T[fNXI9Z4ELR(
^UM/LI]#KV&.AO?TJ#@NT^aNCN^&#Xc\:T4C>[?E#:8<-?cbNICG&/W3.g5\&g>[
@@(M7+W#P+gR=88ObfQJK1A_@d7.Ug5ZDVM;/dbRH9Z42[0ZI@G^-3>C7dbV9EgI
,75TMMaHWT4MdI7>ZW^F6@fYb;FKB#TQR]#@6R\<:AU[F=6+8gBE43=T2,<N&[+<
9D.3W,#f[7)4&3-^2L-LQ(K#&#(eWfP6)4SSF[@HVJ7cB?MHdB#_XABXFSWVI6TL
I)2)aUBaB0O)V<E]GW_dMG4.fMXXWO:GF&T+0DJJ\,8L?A2B#_J1[#UBNEBL;PKd
7OL=VULVJST#SNBd1G:?.Se&[PM+g])ZB0#BCAg3L[?0.c(TM0H4?+I:H/#BCR_d
?@cf<+4BSd27BPd0&Y9G6N>6+Q,ZA;LQbVQ.4bDD=f;E^,29d;12468e?K)57=^c
Yg]:Ae<)bOPRg4BQ-fUeK=,\I)RKA:P:)&Q&F0Q_?AJ/9e=#IZQf,-&2G)6KU_g1
)UXH^]^d)C(01d#^cb]++;P8QfgSE>LFT0&6KWQ1:7U^4(4aW8Jf#1ZDGGJJ]PZ]
Jg6b4a73^g)RRH&[X2;H-;:]CVXeB8/7IB#RN,8c[1B:SD(S+cf[&f\ZaI.@gCDd
K)SAWMES4C0<b_4K.&@eUe;BJLgZNZ]+IMge+SEAF.U105FIGcA/-Y;@]LLg_RUP
M2V\<2J-cYXA&A)RW.O\.FHE^AZWg,>VYU//EO.U<X4^bQ7>c/cJTNeGLb?9A]JL
IQb->T2U0Pc^dfVG7+eU9F_FMM&//9O1/KOa4@:Z21b1B2b6g7)FQH4I7^3f-K+P
,A0<FC5aAH#dW-?X1DbW6CL9I,)f96[/C25+AdT=;VRYB_W<e977553<+P3XPU^@
UK]9V/&YIQGJNQ[@>=d7G4@;)6:,dM9;eJ\UGP3ZH,9V]OFfJ6NcIb2&(L[.VIQ=
^N-\GQY/&P64T\Z65@9;;,2\?.;^O#e2]2JD#aA+@9c?81IZ_UcYW@O:&5/R>H/>
IXR&Q_(G^6GG(<(&\Bb4T#QYKM)X82-(A-S3a^.,S@F,01@?96H+SW2I6#G&GB5_
g@5#[GYH.H6_2JQ?cbDX@@G,T)>4R<RZG5RCDF@P#)Yb+A,:d@SHCOg<M\6=2->I
F@I[&.+KTQ3b?<7?BKeLWCCS,R#;&d/MB5V\^K\069Sc+VKbaY8=F^@\+>X>b]C4
)1RaAR=bLg+EK_CB6[0S5R\Agg]]a@\+MKG=Tf<)N(M1R.][+7<cLFK6N<C8V^/<
3dI.OWCTYANA]14/Q)/__O5Q6fJFDZZ.#=LSgY0-=(PAD#VI]>L&I]f/L0)LS+bE
I+W&+;:;a_CS1@R60TH\UMOdGQUYM?[)8LG+aW99?e<1U._@MA@C8,=c\T1d6MH@
B8)THc;]U=A^TSC)1(2/Lb<e]I^@B_=((J/AMT2gaZWI(#^QMg>JR#b_8Y03(UEZ
3ZK@eg1C6[-5Yc9LU.TY?_3PAEH\2bS^+;3cM:c&H=EB02M34;;YYe@O)T5[d2/g
.=.1]XUSR=(9TF>T&Sa1AaWSGV;P5P_c,63:27;Ze]e^T9LV2_3Q>AK-4Z#=2c:F
4(+QFW&d+]=V(4XdV8Kb3C4UMDB.V#8C=UZRYgKLDe^=gNMS[:J[38Md\N<&M^@9
62R:DT0212([@dPY340@P?U+MZ7NP3_VJC.(0B]LgBCF\V7S2S&:a-2DZQQ0+>@&
(.>9189E4/:O,?5)Ag;,EMAM<>^KQ,TM4Ie4@c^Ea[ODSGZPX2]-;_AJ:B>59fgH
0DN2^&a-A\0e]F^>T;GDT0DA&K#34BHR5MDbE]JdE+eKdC#g#6.8BL_><-UVH,0I
aJDG);FKU..^d)=@E97,,Kfd-64GWD5Le?aeG>-V]T+Q.FeGd]?:(MM/<,(O<VDP
HT@.NGG8-]8S-V<UQ#(:TC5M?HZ/Q^9&fAOfJJM>-G>6^b7g4&-()Dc\OSJ;<9]#
&DL-?X=b;gXFgTf4M@].5.6gf6,NX89;^c5_>\)2SQc1Ef0D.f1,5gO[fWc@^^C.
6&IbeH2=J,LIf/1#[[#UU<]:93N5g#&U;@Y@)S3?JC/V)GQ(+VC-gVNJ4LCBQX4P
9_B.X/HPQVR@d1=?99:;N2):HO^/42JF5f-8K>K1B01W@()@cd?<O-JL+=ec]1UO
f]G76)_CQG0\-&RU>.ROU9fES2-_YOG&3J2;a+-994CYI=)G?JH83a3(d9W;PTVF
F:WU@GNHQ2M4SJ@ag)82IUO<41Z5OZ]AZ/,5ff.Y74O(2[D1KPC6UOZS\I9]#?2Y
ZBW\#S)^eF#+ZK-:LH.IMBL;;+S)78;fP\F&)C,;>OU>QJfZga3.SSYe(EWJU_8(
^SCW;63O7(\Ja^d]NB:R&EBBYO?HED\7H_?]P@18b30J<4LA_3.5VZ_CXL/fBAJ,
fTb]UGC0AV5fMLI@:)7,R3Qbb1J..;5DB]Z],)B.+DV6YYd&d2d6TZ.]<U<^.A>8
NTNe)UR\5W.)g#Hf?6^a4J=P.0);NOBWD)Vb(b[[KOdRB-.ODUe8(CLH;)(-QOHc
DeYe86ZR\=OdUdWOG4?fLD&006VDPfA3X_@ES[5/cVe>Ec88?=U&JT)3X=:PXG-K
VeAfL4^@M+aQE&PUG9;\I_]N\+DP8>\WNC50<R^SQgZE6?D6T>>cZ7V@d&Ee7\51
W53aA]+Z+A:J5EHF+.;]/<NV0W_QB+gZGRFN]SF659dDT?T)&+_XF1>VWf,T2cK^
3g=]Me=NBZDT;UAQ>X>)(LB8XQ[J,+[]6g\(KR7^ES]DMe?WfLBE6UHeG)WNW@WE
#8K4d>?8e49:RSL2LFD<_YHX>04WM/ZNXIJ6I?#J)49.Dc+F>[RVE6(H-gO81GB]
WH=G>-@YJ<@)VT^[X:D1/]]QKIKY23HGS;OV;+?Q=7(8AgTU>+1-=DEd\L2D94b0
\B<0fZ9&[@0N?A/5bb(RII,f3W=JZ/+JdaCB?\FIM2[>#I@7&;@K1+cP-86PTVLY
Q,(TM3Y^I/\4BfX]:7.+5fg;cFf5?OZD?U8_[fZOX0K3F<7=3AYR5K7:gJd+8NNY
a4(JK]G-,g4:I6.4#fXU)_d77QRYF#OR=TN>JP@S47HadI[\eG,a;M520S&H6799
73+F7R\D]8TXYSOAXdV3N2.N1LcHbKNOaP8ffLF+#4#L>SDYHI;611^7P6dd.f3E
4\Q6\&BK89+&Q^RD7-OebfJ:P<;>Q.75@M)_W.3G-a^[BGLd?:Z:\(88QXJ0.FT9
NB?:BUc2_<>34=gd)1.>d4[6eD7F:X_/.0NO?0>8]CXGf>L&8\<c[4:acJ)-I=/9
ebJ5M[/Q-F.B]6@N3&ZE<d8^CO9>7Z#ffM@VD^5CBeePe^VGZQg?N?@eHNG5#F]@
DP0dHG#NECOM9BO:;RI.I[U)F-Z[0aI2/V3f9<K1S/_df7&AKS2B[,S_,eXT41Pf
NV&PD9)J?/#QY7CZ\[VBXf)\7[Qc\N^_0#(cJ.FP5[>A4U;6V<D[F^&B^8-KYb/5
b=&IK0;28SZ=HC[J2]E0=,D@3#JSC2@ZE^A72_D<J0b=.bg6+>UAL,IL4_.T]1#J
]YZLW7_L8X[THCOWeTG.>/?F#A>aYGZUW9400:L1]RU:(^TK-(@VD9CgOQP+2>WA
IA0c38YT@#R5KX\^M\[dZM2T].?J34_fQe.d0U=\O6N++Y,J@F6.;?6RL-5HfKfZ
8b96S^gG7?WYW3_bPc+/d^LZL8QUZ=9Y?>F=;CEID8eN\#/)P>aP].RMMQ.KIY45
.RL07]?(HMUcRY3-]bF.R,SS+&:&4O&23<)A(K\F/-8f\>a^2\V/:-EEF5d^BCOe
M05@6@?JDM@#=EDJdT3L9EIbGOY2IQ[,e<_)4WR?E#H8+/5WG2O+=G1c[Cb.LP&O
Kc05]T7dBBQ\PIEEK72WXb?SIK-[3WcWbAX34:;G&SU1#0.L-Y06VLP^5R#0/(.G
8f\eI>>B7g&YD-C]EYBXGWN@:Z2O2916c<\F#a7CB&7PcSJ&#0[cX2f4]@G)aZbe
+-75T9\8VJ5:@]Z5cW>Q0f>,4<e[D\gU,FP7K,J1FJ7YFG8D->IHOYUSZ5F/PZ0)
:-0_LWIGBD@Lc6I[<57M&Y[e:U.;.NV<:C7@[\LPcH7Y+Of.EdHFd\,<c_;2)FW9
>;)-C-]CaU@f+5gX2U7;ZB]+WB]H8S5SMEKU@RA#43=Q>#/Y2HW6GZbN9\WWK/5?
ZCLU)<daJ.F]PYZe-]=_Z2]]36ZK_/_8cR[#ScE+a]FBf7,7S1QZSBc?NW@B1K13
4U/dIYfZF@M8K22KQ7CG9NZM[E9a9fNaQVH.=,O8X4N[<SRfZZ7@>=@XO]]K9S0T
I]1B/;?a&GMCM0YfF_bN/@6GY8AT7g0)(UNYB6])A8&Td9DGLL#=6(E;MABAF/\Z
W.XFeLM@R7;RT-]XTJQ1Y9XB>&7gE+W9_SZ3gCW5R>.0RT?X8g.,:RTF])K7->/7
X[X487+4[YfR<?+^X#]Y/F_>eZCe3c6O5I<MVV7cY/B,eBX>/4L7NY&]78RZd@]3
Re#^Z518=VfTO0f+CYNIg^ObV[V04cE3a&O;,S-ac#PG(QJ4B.S=TF0L=<]Hc7&>
OD;4H_cYZ>D8ZeCGS7ZZ6S,M;.PZ#_?):1I1c09Wg1cY9fef=J/K=/T)Sg.cSX35
.DR@71Ed_EQ^<H\[X3@bV=VSBNWR+IW=O&PXJOaNWMT/(RT0gU\g@[3FbKW8,[A)
\59:d>b#GeT9&&-e+FaJ9]8FJ,0=S\^e(c+EY4-ScYe<?>;ER-EI;d\W(JG1B/dX
8bKO_aVYPQ3a.]<eIJXTLSB[FH-7J#DCT<b,:SW)W;\0K_NLB[,T+2[H=fE)\9VS
#^fTM2N^W_^R@39GS5@=cWW<;54]W?9OUSEV6?(;BR^8&:7_fdR.ZgM:;L[-aV6a
eJZc0W18C>2a\0?P7BJ]/Z37;Ff804eWJ:-SeZ7GC39^([BTIT6=c<GBC.2>92X4
0<J7RM(<IQERS^JEQ&)=(E-;]4aQ+L?W+G<dN.b/&8[/#9bZ[D2d6HL&:9(I7.E-
QU.KO]?f/-]IEK(ReUTRT]4aHC[V-B9>D:LOST1O-117T29[T[30;YGF.cQ2JD]b
QW)7:LC(;HaAB:7WH:?1<VD(TVZ3K?Y&G\\PdQYg8N\AXSD\L3E>He[)=#;^:2)2
UN53Y#FX01cKCC#N#d)F.A<@&5gR5Y>&NQQ+_f9[XXL9Mdfc)e.Sf;0-\?fC29^b
O\160KRB9MXM4;<K=b_D5:eEIAXN2FTI;KY@@K-P;3^[#gM>PFRf9XTYNZfGFU9@
I6gFL063[#R-_eXc26;f81Y\((cL#NV_N,c3)B2?(AUQ@E)96O<6\d7IWDACUL6F
Y?B#Ha\3OD4VNP@8::#Q6_.+OHTR+<\1N\3U?S^N@fcYZeO?BSbK=.<>YFS;_/dZ
+a(]J])_^ccgXX)4LQbJW@81+B^EKc@70LO]BU4\RIA5_,@?WF=b\PGdb=fGK(Ff
2SMQ<WPa\&bXJ?XBI&1\9[@RTf8+7V<g2gT7T<dIZ5^]1GF[J<54Y??,eE)>eSe(
>8BWQ_efVfU5HfKP0aZH.<TTQQM[Z,Y#0HXR>X[+(QgaH\CT[,K<91#c/Vf5O#FQ
06EfA?IgP6g:Hc&??-:);G79bE&7K+,5?:,QTH+)]IIN23\V(<NY9/S^=Nbc46d^
AL7@gd=715,OIG&VHFC5]+bJ\)\V);_e(<H@Z&Sff2&O&NC=;H#)<Ba<9H12P,/=
d0F+N,e@KOJ71M35K(X.8,?Q3]X/12K6+@QaGJ95DGd8M.#\1aRTd;E7VY3XLb6H
P/@DQE@:[>a7A=bL?^WL-=IR:E2?MV+B@L8MXWK<<8PJTUG51Jb0a@C_KdXJ@=UM
QJQH7Z,6YS&/DCEOB1H>)5gYN:=YS[WE^G-(0fB&,H\9T=/K[&bUBKUb,^ZN5^J<
SLU#<K[P/ID:4C[UP]RP,]WL(8#RU^\HX_\,E9:;8H[,4b3[RF=C/UdZ.IINCJf,
]UEU:fRHZI,#&+-OU[b^/ea;]4E<?^5<TdBSKC[._Ze:-Qd]2Qd=PI=fZ)J2K6)3
YJ6KND^HG@=&,P?eNFHIP-<&:SI7>ANR8J[_\\7YDf[S-XBX6ZX)Q::82&Sb@B-H
f3O25XH+X0V,5S@ag8KP9faM6IAS9+<A9SA<SR>I67T3SV\Q^O27XE]\WQ@A/.^T
#HS0;_^>Yg[RIDF^-T-216d4cXXd,OJSME\NALg/HgOE<Vcaf93ad0b<J9UD=BYH
cMWE49NUC1\LC3?HaB2)EeSX@e=TZX:_Kg[cB<YU2YTF:#=2>K>FA)YONF;cJOL1
#a4RQ9A7EIYGH9FJ(SC0;:3;WdH./UU>e3.R)?;)1dUIU]M?0IZ1]7XX&5.TWZ=]
RMfGgW.?ddKNP3NNaPC>C<QYf[..(0].bcY>)dg-TB<C0W@\-QI,bJ9_D-U,,QKR
^3+MaZ72<6c/:+(aQ@15K+Gb)gS[LQF-X1RKU(U@EJ8/9=Y]2YbIBde(M]K1),EM
f\+^+),.cNe,>=CUg&^gM7M&58cHPN1\LJYZ.f>;1b:X2N.H;P@WF@\B[U.AX\Jc
U,g?,9;IS+)8#E-RC@[M6ZN:Y0C.L33+>>OAI24&</6S.P;J;:)TU&XTcNX,\3)C
E\R(J>4&C=)N/YPC6BAKeW7DWFD<Kc/eG8gd[0.,/?RGTMW7d=d[.]@bbR/ET^<&
(RAYc-=A^[FF1<Ia]9<eEC\?U7;U9W@T[#WMYW<^>6@)B<:S^O8R:f\HEO3\/5\^
UJB)J,N&a,I^M>#(NI2Og^^/CcDa]OP^bdgQH)X^6XRI4Q\E.E=PgK06(dYTZQgO
Vb?8.3:48fO^<ES)M9Z6eg-=L3d_UEVcEC==\I13@6,8;.ObD\X;7XRd##/e#=((
QOKQ-_Yb\Y23@7RHEL+#b#.RT[6K^,=(U\#,aS_]7;bVSL9:4TD67eW8(e/#+RYR
4,_12&:b^eXQ9N4Ye7H2:(J/#g^g]55<J)>;3M//SKe)H^:DY_;2Z\FO6KJ(G5=f
\ADURDR]P]96,ZOB2-0RF/DID@V;eVIdS=9^)BB:E;OEZ1QB8SKRDaT8P4IU2;)I
]GcgYN.TG]0G&7B4XTO0<5A:#@Wd-C?HDCH0=BCARGFA<59;;ZO^=^&Y+VCY(;)K
0O1Q9,,,f(AZ2+N3?P(?\D8R[18V1.QFe6Y,TE2L^RTgP\g6T4[E.Z\H+-#-05XQ
0<W-C?#&X(M()[RX)LN3YN]80c_5[]\8#DcBaD@7<bF+EeKTX89cc^N1QTd4;:_V
cd2@866\&B2aG>I-,0K45AYM:ZAX+C?Q=eIbdYge\Dd</&+[[XAeGgL+6b@7S=Nd
b;Zc/MX/5?<BJ<?&-Z?[.TeV6R:BMcGVd:Ue--ZKde;0U16S):HGb6TRU/)fHR<D
SfSO+QaKAN(V5GCUS+S2,cFcN-ODPJ-2QV>g@?G);,7Pa#3KgDeY_f0/FPZ;gGfH
]?V49O2&U((JMJJf&_)aW+8MNeQXPE+H,]LEE;LbL8\Z4,1YIQY.@1YL;QI+W,Zd
22WPLZQHHYb.+7eD+C42;Ff<W\KHc[@cU_deB/.MX4Z(R-L[ELeSOW)K;WE_0UD7
AL)2&5,-P_R-EA&=6E#^,0@B]-BW4F\3TBRZeLOMD_0DN_+MS[SF/:EV65VOWcIT
C=+4Rd@:bY[KL+(#R[<BWfaH)P2eHP5W&(6+gbWHF:U,:7(:aV,0e2V=DOaM#HgE
;4<Bf,+2G7.aC+4\V/KODC/YC-@],a\&72:KI\M4XAg)S00G;3,?,P<:FT/2>Ke/
9F0Z^Cb6C]3AY0@<>9R<:+M&W#F3Cge\T?G&P1BJ-^/Y3BA)1+dUER03f2UG:bR_
DXC_<IREX:85<S9(9FU\6^0B)\&0Q,d:7^GLKR5S(a#OGEL\(@J<84?eJG599C6d
3F#_c9^1V7C-OcK+G8N627[Ad^;89B@(LH7XBPGPANU1<2/8[Ng6BTH/4.<bY@=a
4Vg[QEZeEA/JMbOR,TJ3=KBg;NA8?;L5EX=f8:dS:dG#&&4OZ&UW[cMV/^/8Y[3X
Se:(F7D8)YUCENeNe;9WDdEL=4QL3@bde(_4T.cd9aSb/LggI4CTGJ-<>6cZAH75
N<[]3U)+[?B-Q2_Of[\9XJ7-TYWIEM@1,RGZ,](QS7?A5TNL>2LNW/g2aAc@CR;M
)\.1\7@0BDYBfEP+(<)I5L#8FG?-(c:6c-a(5:9cbW\]&J)(F+I.6eU6P^8/-\V:
7=)GWDAb33E/&8=T0?.R[bfC?2:J([/,9NcCG5;.@7gJQ.0@4PfON77.118AH#)2
E2PC1Z=4a.O#=@MU2DP;9XcaPP<)O(HEcUNg@g\1(6)GB5&1^cX8NM7We9]=ZN<+
(1?B#LF#5Nc?6ZB[^cQ-)OZ/EO?];F:;b;_a,YE((L8T]8.E>/C.2?PTP.TY4146
?PC2WUZQ7M4(F)J5D[XK:W@F0:14=dQ?>MRgKdgU7&7_DHPDY#SM/Gd(.(X_.<JN
X31^90+CS3C@P.=U(Qd@43@f.GOV;8JX7C\Zd=0WHEK2/1)[#9.6UI\IUfRK>[,J
=<-a)M1]&EM=1\6JT23OJ18.I>W1\GgAN4GQ;,_[He6[-3RC3N?.@Q,SW3MI:c@H
&-U9eA_3]g.;Y;0>=;#,8G8eD1,:]Vc5-WScB(/#e25a)b\T)>Z1+P#\)H,B7338
g^[7]55QC-21&<TQNBJR/e7Se(KeY_2M]be[3f9X9INd/CZ[,7<8Se((@TVPff3.
AbFHML^BM<@,ZJE8W8O-^E3KYVMUfb;caL[&Q8)dO6/1L,/g5,c95@<-<XS+2O:,
dD8BC#P@/V?&_(])=0.ZH9C<3OE=8L5T_T1:;^ZBOMQ([Oe1Nf;_23#=I6S7fZ2g
.IXdE0/A@RI2SOA;9(HES6b7R.[YW&-/G3NVC,adZ#JNTURA3V1c)[FZX09(0e<X
[?Z7,W^T_7Ec4=P+6]-<HN^b+4S?>SYUA2OJ8@0/N_NA;43H]N2#ZDT7]>:82F;Z
M9Bc9Of=0Ode2BHB<FcI<8:1;NNB252:.Ab9]ZFL,)=,SH&aEAUQ3;PD)c[8Y1T,
85=8gVR>I<;/XRHE2(+9Wc8W_bI#;VB?XSSXd7N4_77TW/?,OD\#6<9RcEC7_R#-
c_.F?g(>++a8_gQTIYYI13(\U.CD<DGU1I/WN-^#-(Y91KeRH^R]TZ;YIL;>;B[=
-Y]O=)X(RA)4SZa-QT?C>\KIF._^9-P2;NCJ3He2[4[0:C<OZ:&>8-d-2GUSV<?f
ZaG+8U26c6IGI:aL,:9[4Z@aG<c@0:.@OCBg?MUQ)T-K;SNLbZd&SeHWJ@.V-6?b
=#0&?17d1;#e#;\PF_dZOA/C7YWM0)Q32283Q&KcW4eB#88N@^(92?0.LTL)f(S5
DB#O2[f8L2<TOdcWRH;a6C]V3<,I.ZV1)AY8?&ZW2bI0M_Yag-N-c:HK@Y1EYLN5
^K_)T+C:Yac5O>&C+7&^+\W[ab:8PDRS[7?5Yf)gVJ&.A@>5JLCgMDd@c+PBC&.8
M^g3&X?=Y^F)>.<W;;2Gd>Q:dTQQD;>G_^Fb<Y]H_H)6361\TJFC@E[b[Qb1fR98
4(),L;AD8?D:,OG]8R]KV_@f>94_WcKeA1S9b527>Xf>W^eEUQY5c80<E<d.1<JB
TN<T:6<a.>g[ed?Ta-JEe_D/MORb67V)Ud_Kd4P^WGS=-1)A[[3g,Q>agR?HcN/4
^I_E(Z]H6M><O0V#@(7)S9CVF)FHRZDA=#<?G6[EH>dCG[<8I\d\L3O&PAM[^Y5U
:J-2Bb)GK_P3)gR4<YB]@acUbeU&5ZINUMCH:-eb@Z_]9</6+D[5SZ+VY,H@aD/&
GC;dQdA(e.7I54=UJd=b3a)#\R:&E@HQZX6OC9ce.?73[CbDfd)OG/]6+)9LV-ZT
Z-\e#>HH70&IE9X;>.fZ_PaGOOf]CZ6b?LO@W8_Dg,NSf(OSK.M:Fa]NWU@AY2;H
9g)@KFL=P;M#NH1-&-2C:NJ^;:N:.#efBRH:<(.#<[_bX:GC3b,V&BRNLU,):^R(
2\adZU<gC&(eOES_=0\0R=I+A(cfGaA4>/P9c;@(FROW6\DUe78^e=8\@d7QGL_4
Eg=g_\EWUP4VHKC^C7D2f8F#VJA=4>.8;J1>b.:[)a#Gg<L<8MK1TN/QgNYLP99+
4]De.0\;_Pf=^Vc..M(KfJ;<Q47PA^)V2X78A:@9]Q11\-\^C_6JPeIPO14#3LBG
_TW1(H[d8_W.@_.cD/7dT)C[9^1^FD5^]XgYOM.XXTYS([JbeA&H[2NAR8S,JF&T
0FWT,1^,YL)#K6DNPE_O]a-NMK>7[7f\X;f(Y0=INQ\9QH+G<LZNA@S>6C&Od<4b
7LKDHf^/c)[VY=L2ED\Z=\R/,8GcZa9UJ.O>B_fB[@]VZE(6eDUTg3LK<VFBF<e/
9Pf.(,?V/6.a,Q?_9Z?U4P>#A4L#FU=E:fL,+N].4#W\af<7^XKKS(\N;2I<X0)A
1G0O8Q4#B3<c_9>XXCa#,/Q<57E?=_Ug72:KEe#@H\_#aNEG/Oeg0SBA[gO<=XaA
2fXEG+a/3XIb0SR&Pf>eA1dBOe_08[OPFX+Y^NYC4Y5Od@[6=877XQ;#dA2JN\/?
aP?.2BbYGN<\<Z1b+XQG)UY)QDY++eTN+NDBI4X[OX]f0EYTN?J4LcAaKF8dG7F#
X1#_J;7@CWRTGTQB7&./:<IfIL5K9)K-Y6S=8M&C67X1D7@[0XJR-HLUB0@R1P:f
d2ceVY1CM?KX7#b4_Y#1S=7<dHC8Rd+;B45>^([M+U<50^6)dP;UMAS?[1>?#g0I
7ac/E9VQ,_VPOFK]DaXfg#bQY3:D03gE3Y3Od+Bd0Q4?g_SL(U_d#=;-M&6Gef6&
0^EZF2FL[>7SC8[6fIJ>S=/13M<L9]]2,-WOS(1EQ2V3&\U&06MXY67?7E?IPJI:
I0@)a.0e^VC1_ce1([O7HUYT2(c+E]RA[gb;RFNL@?:a1LFT](^QKTI_X\=/3b^0
C&VTJWO+3g#&_VD4;6:a\MON[Q#F?JZADaDD17<2];egX/>9Vc,7P@@bV#+XPBJ\
9/_c+<(OdUCa]DP]BKY9D4UBV[8_Ld22M(-N^XgCJM:>2&R&Vc^^dOe)bW^D;4-R
8baW,bD);P&Y(THLYV#Eed/@MO7;0e?eA>]eXW<<bKg/R_Z3_gF+W85(A(E;EBI_
<gYX+egB,5R?)7N>9HBc8[3&.?dc:(?=fWZ7g&]_[A?,F;N(C7G4>]):2.;T0TBZ
UX\/48IEC02;UC6LY(#_0)b7,W:bCJ+PVYa=dVe<<3FOcR>BPJBS@\GVRYO2a+SG
e8<W^)cRF?V^<\6WBJWI(?eWP(=#>#ba-9\\5F/L.,/VPV2c(Og9+,):d^XRR[)G
D&-ScZ2)MIA<aJ(e>dB>e00QK.V4TCS/9Z[c_]dA,T,+O]aSG(PVf8WF/;65:).2
NA=7HN?\8;V.)61T5PM\V.C/98(9Z]#@aR9Z_bA#]B4GIgDb)f5[Bb;XMd>])NAU
WM,2:cFL23HXIW.L0ERJ7RSCR+=AR>;MR0R<e47?\W3[F4WVHJgN7e[X:Pg:-7LF
Z^2;cNL4:0B,;&U1P[1ZY7QR51fK9H>3XT4)?RKNfU.b;+gV#UJ-:F[9@<CGEK.f
Q<dade&J3=Y++VXG\1Mb4AC[<LaZ&WOFJEJ(fWbe_F,0)OGE4IdQ+NI@3,M<UF;O
eFQQGJXH[<fGIb-dNBY7^Ic2/>V90eOIdGW,X35SHQ[,XFT:;>P1ZHcJB]63a165
PNGW)6f7-[I,[AN;TZ>RC)D\_>E)T+UYM4@5+H>;Ie0T0Z.(7K07FCa6^4=5Q?/&
(E3C.D5f.8SOcZ<\L<T1CSR-<KD<QDO61[X(PK>-,)&2L)L#;V4gI0,1#QbT\<<M
B.O2IS@M6,P8L1JZD6@I-b9V#4@..H.3<e82dZE37RUCR5UH.gbB.7a^LcV?RcJ^
#eKbH#1+_T\+adS&\aWP@8#@F+6@;TTeDIA9.,MRaSC:)>UY4ZRO1:R_@Rcc4D3B
(7(+2WVV8XO4=@VG1OTEFX6a6A[,\<=YO^;UD:][LX::;(c6f)NM4BAS-=NG<#W0
+26W/2UBVD7DWP4;_?AZT^9Zg))T>1Rb@D=6ZO=[f9A5-8#P,Z/^Aa#CE763]+,E
=CABeZO22Wd8/B8(DU8-LeMCJU]UcU+0cDHfC)J<,(=Y&)T72(V?Q&<1DD6]9>4#
E-JD7B4(c?BO<g,J)-ce)VU]+1ZA_I8)60)a,D]bM&YUBO&^e[?068P]f2PW<;e,
90Ea8aa45g=Ob:Db5]R3d)O/\P([E)]Fc@+^JJ&1bfM4WLQ-_5eK.Ge-+7:7NEYW
)FcY:RCaQg6]bcB<dE9Y@&a232C@@@D:,bDQScV@QWLe]L8,SU7]V-VH1WX>c\U9
-gd1>gNIO=g8+dbPTB0]RXL,;f:V.d,3PZ?+;-Y)=:g8XF#KFF=2N_D4/cdG&U^Q
M1:)@@V:B0@Y^4fJA7fCQe4+Ag7cf_)97&#YN1TZ?Zg=O&6^VQ;X;)JD_4IN(]G^
WX7cPI.87]_aTKUHE7Dg>UWX<_8L(5HY+FXQ#5(W+e2V8=4];,R;7WG<,U3#SgE=
M7f\;50^TfC3_@D>J-H^0I>Sd]QdH5E?B:,#A(+/;c(8NRQF0P;e,Ve]MG0Z4HEd
V4?6&=;cF9DSBCdECA4U_HWW89JUX.G;A3T[ML>4+3e5>)gR]&T3AE5K=8K#_LO>
D52#V-Q#YY)3NcEU@_=IJK4ASg)aG9AN-WIG\/BECE51P9HHU=I_EM+[Ige/YAf)
5K>VCA<3&c^aYAFY:71KX>]2018FZ/a.>+KKg4T7G]=[Ja2,@7^C\&J36G#PIJ1#
/VRI]9D8/fM3gJ1cN.U?.Q3N4cBI#Ag_c7d+;gKP&BD:dSS\?S:SB8P4T=XS_-ZJ
J5)aM0#.;[D)@M;0E5OT1]bG-93Sd;NZJG:55XL1DJ;RN6S(D+G@,Q_DZU19;YB,
<(0FVF9C_GG&cLR.7[[G&LU>QDc7-]:FIK59M_/#SK-L^bRRWK0NA/e77OY,BYaG
c7<?LYc=\a[BXUa&,CbI;\/1Q()^CLTWG/T7.F-_F5ee:?\a.SP[2Lc?ADE)PIdR
e>4aZ:e._JFE.2U+b86O_\FVQ=.8c\U]F?(UEYa;DfAM0.>ZIeP&eA6#5OcT[c5H
V=6:=]3;,BC-=c_SR_-H@+\ePAQ;Wc2E&ZSPO_&=4^4Y_AX.+0RRg_,68FIS:#bQ
#H_?0MBfe_8]@HgR9TMJ:X\<9D?W+NZ<)H\0H-]^ca9CeI63BVL5LHAY=N94D_UI
SK>7DW5N>H14#.<=DJC?)T,,(ZA::P-J5DVO7^.U](/2Z+U)f).E.:=V-+7&g=B<
LG?TJ..O-K::XTY=KXTG@XOK8E<0Q>2#7MJ?>876@YOB7G7e6/HS0JMC._^MTf7#
5(_P/^P=M<IHbS=Wb;<2C>3OEWO)APG&8=M)V:TUPHRbIb6Ha;O;(=^:bHf9R&+S
AMf822^^(0T4HI6+fg)B]DVR2P(Q:dDACdDKggU<.(fHL&9]ILW(&c.#D4MUe_/0
bQ,NZd-g=^9)_(-Ycc]^#.M-BJ1eQ/#0&YA:^>4:FITQQ:?YZ<VERJeeTD;&9D+O
B6S<UV8^d_HX14?5=I,JfN(Q5G.(1\?+F(_6RL.]gYde8e06H=[84XLWJ3XY&CK@
GZLZPf5W_e3fU(HYXOc77R5HYA<LW>_]?>>&EOd7GXTYRBEZYUcFUGD2)2O8[[)F
>L<1(4c,L8SC/2BKHfQRENQFd)5B@0#P.,A.O2O[\6GQd6PUV=c_5L5UG2IW1QX<
L(F#E]TN1-]Ba&:].]2b(YE6+YLf6KS?QLQEZf]+\5^gEA-bCXYJ1986L]/:^DAU
QA9O_P0MTa,H?dJ/C(,:L>^JZ76<A9E/Y7gH9ODNRA/C^7>BD4.^@8Gf4T]#:::0
,e3c->AAIRHf&Sd+@HCAP,Zb2TEAS4Q<[#S4P\0<]L+7X-D39a+[_Q&MU>:50)QG
<H_EH&e-+3f5BQ=2N<TP;\gC0;P+J6=>UZA>M.[EFLT0:SDGIfRa.QKc?VPK6\^T
WP@b;dc.)F71K)f3EYA=RDSCIPd_EbTP[(=RQ)3+3<M8Hb\9cQ&C8T-Ab3TLdUFF
@T#+.-4b1^O&42JJbHN1;A<>9e^RE,cX2(Z/]0/FR[>5[Y)_V&U/M>L1][J,:91#
8F.:XR[B3=THJBVS))F_KCBcbE>F6FI6Z&BV=#J26VP-;0PBM>#PR3)9T+,>c9<S
8+PU\1:BE8Od[5F(UNFSPON>/e_dW+08&#d7U9cVP;J,^bebcaS@DQKF[Ea)+0LG
^S4CR0&_VDGP>/LNH(cR+@[W47K,K#.BcECaX\Db^P4f2@X2\\4E4W(M_2G07SHf
CXQ:4,Nf/<IKKC^O9dc#DAdS?CY-FCAKaTAaAIHX]SUPbWg8JKMUD1cF=<#F;+?A
d,_-a3:FWL)9W=P,I.G1(H6@F\Zb,]/WS#=cSdL8b9^3eT=/\Z:)4Pce[.S^1CeB
DT]_cN;^TML]B;.T(>49a30:f_QXE&^49U#7gf<a]@#g;9Q&VfP9CcOI,e;Rg&YM
BWW(c<Va0A@(V5b#-FXO5N9[06B?Z7TYIAV.EMcL+&I6RE(4RN6O@K3H[F_6_H7]
e.EgTaOc6CEDQbIH7\#BDK/P2>ZARUP=6.NWCP^_Aa_JeW?T]_)Fa4;K+GM/Z=RZ
a:#CVLSU6<),S=#VD1;\L:fBNL\QA#&/F@]>]afb19]?\fR#04^E[DQ\=O0d><QR
#BOa-@Q^[gWbIAFg;WX/C3ZMF,=\IE0(\+,M/8]:Df007_ULEM]1Y:AS8H5N3C?[
9\?X1+.BeMc;BLFR_H:4U@-?Eg38QBKc;>[d>X>Zd/2L[<Q7]K))c@J.3:M^W]_P
TLgb,+R3C_1=H@S3[2)@Sa#H#6]>gZ\-5J+MYG(U8N+;9B[F?@J+/-gHO6U&=E&,
9]eWCE>_gEOcN7I)@#,dSLC2fT;4KHYF83^B6aI<VH0F=D4R7IKH^9?gc5F18/AO
_aI>NT/GC^P>DN,4Y_?(ZE[S0?W#,7K),b(XJL:B>+MH24=03baOVbL=-O5)d]Aa
\[YT<8[f2VNDe]Q?+?eN14gJd+,BS)@U/ZWY_WA0b#C58e5dMBKBB]PZZ]<CQUO8
T\])dIC3\N.WcYTKO<;AMeG.b)YJ-NG(QVNVBVT^=R=Z\[<7OSB,G]cA:/2.]UC1
717TLJV@6<?\N8;0SUg_d,5JIJf^)gcM;.?SZV1B4X/#c[FbfAXC6SaA)RdXNCT@
]1QZ34GZ[]G\PPR]&adG7ESfe[Ga&MJQ<3c)2/Rc@?XJ;&&_6X3#B[TFKfa@FA-/
[[cR,_;8<g;X4LOfC3.DCEB,L=/J-Egf,^22&FQ6g#MZM9^31S+C6ZAD3]I9LN)Y
^Q?/_I-ORCda5(+=W8S-U_2@Tg@_-DKS9AL(U8)>_NTLKKF&F_[FBYMV\J9.^&]/
_e86Fe@ZWb^3BD^ZV#[^H5LZ+FgST&Ef=P<Q65^9+8;SCB_,\E-9EcUTH:F=IE2c
2S0Ac,7/./S55T]4V01^&^BLP7.+K,+_.C>\d409/-O+/g#FUAWB]G,>\I00M&<M
WV?LdI4KY86YW-W26-)5TDQ1N.aA+DKN?N;29^0(eGHOM.XSK;>Z#gV+b13_bD)S
FbP79T>;R<KNW^REbOb7SX+I?6;T\VQ2Z(H]Ua<#[AcR.UB3aN--AOSYA[TU(Y;F
3ggf/N+ZKaRF(+ALC2ARE6_AU6_>^X^M7E71A8/?P@_fD?&#d651K?:SLKXc]7_3
GPL69W77QE>aGRY.R#+A@GSM@cYBUR5BW02ML,&AE<QH6RdK2BbCDCg)W&1MJ\J.
b7R>\X)39WIc:8fS&+_QMVZg(+<T(@D9RJ2+W40LHMXCZESL^ZD2#eZ[,[)LDPO(
EMT:I/<U0B(EB)RXNZJT411=7RLMaYH@/_BKZ#(Sfa@DZS).BVf-:40TY8/]Q#CS
.FcOL5&VTK<?PNG(,)3Gg8K;3O>Q8B##XS5UIT1T.4db;&@D.RD^dZ&)Ag1<)U?0
^ANEPA8,E4(e@A#DTXA1KEdf6HGPcd(S1?Xc9#L4@ZO5dG-\SWOA^\2X0H</?4&P
c;Rg7>6E8W,I=?O\]4;RIQ1cDO>.JaZ76<]C#QGb>^BF&;XaCZBO3,.0Hb<FQ@]:
KH.5b5L#T:aI14MgZ2beYf=R+?M+E:a&X2Xcc(.gdbf=NQ+4@CD#[f\e)Af)0F[=
_B;Y\b)^&?>R2;JUd1Z(_T#.C-[:<SHQ,N9RQNOFf20/DB0=,@,90Ha0OB03DOe0
gC>FgaOB9<f-14;A,VX5RH>R11Od3cQ6UgM.@AKU)X-/_LF@#CH0OHdYFIN?4.A,
Rd3F.ME-_NSXeMgN8f94<d[g==P^4gZA##HE5V@V?)HWB8DSd]]cGWP]@RcS0-57
2UTJUINY<3M(d40KJQ6eBcV&5#H&b&XE<^SI<&6TSV@1#J;gPa?B>:,QO^gfM400
R]PTQd.:VGcV8Z.5PRGRYU5.FQ)8d?+_NQGe=/.^VENL(0\&@-#VZ?gc#,LS>gaS
8#EQL7:SEFDK(9W.7BB03SbFfPU4BWO/Cb;CSKM.\/e(5+;W<gg]QD[T26CTI(3M
Fa@g;M:B@Q6;F4O?2=2.)ST7PeYMVOV+E@;[3;0M9(M68R8[-AOY[STM3TYCPdf#
IB]b]>.+^-cE6B)a0B&YC6G:&6@[S^Sd74/)R9Y:QeI\/A,e7cZ>^+5&\-@<K0Bf
J=?8-QMG8JX(R6^KLMSMPHffW2Hb9fc-0Cf4Z3bBf=c8@W5?J@E6MXI/L-07>d-#
6]_T[MU=IUP/5TT3L5-W-/<OH)Ad(4SQ9?9Z(FE:2X)f@XLg+50<RD,./b456dLb
g8JEH5Gg#LXdXLYU0J<-W)8YAea4.b:@]4L5//)3Q5).#f6(g9CK_9^@e5:P8X]T
\,ed2V+BLDL=F<[0>:\J<RUdZ8>aJ\EI#;KV4I9aAB(:VP]@QLJb;#D72YK+g)76
OZ4^=f]??cFOW\JZ.I&PZ;Ya_=9B4<S?dL4JGJU9A7;LFI4N6c>ZL9X0]V-MBBL>
0+GU7\BK)2cU;A#U0K+7RD[E6?eL8S<RdVJ)R&;YO>IEMBR7Y8#&H1N&1<#]Ya6G
7BTRHNRN:c7D.>=<3MUL6,Q_ZVUN95V+SG-DU^@1S^@MeI_a4V7S(>PdZUC8+G/T
C_PXTbBH>NT+aRfGO]1-YEUDT.UJ5Y?9Va58fSASU(]T7OE#X&B[3]fAIbI9/XeP
JH/QA<NQ99g9<H5d//)K[ad8^S[N2#69?+Md_WYV9g;:F;ZGOF&c7I053IU<3PQ#
e9[H0Z+bLaLQ9K72_]00B<K-+OGbcO6;-JK>Xa@S_0Y7,>-L#ASe:]XI_)S)IQ0A
J&RZ&a)U:\57QQ\<>A]@#P.-FYA@fFR@#X6LVc]^a?L#AYZV1HTIVTf\@Q1gSS6X
W#E0Ed-^9S/fbTZTCB&\IWe;C&FGQCcg/?JG?\aJ1KT[@)9MC;5IH#HgLCgXIP,3
X7_eW.5XET\:QAT72-5BVIc):26B8K5RU8?g+Le]IcRY]SERgJP/=fd///=1dK5W
4V?Ib2D5c;E16?=M8,e+Wf_^:QP)U^/(fb3L.^I)JP52-AD6-<GGST)WM&,5M21(
JW12)8;XPCOb;38g43\U1_1H=;A^N<L/Xa&eX;E&+T5>7>aV_A[+.gCL,UVX]e;&
bVYV^:LS^_=E&13K@GI9)M2?eAEea<3@:gKL0NE+,EdOQ:]I@Pae0<+4279g4)P/
Y^O;=PF8e.e7,=&+Vc=:MTR1H>^2fJK?22fZ4a(Df;fcDcYFT/gcV\.LK@)F&dG&
8Y@TH^?Pc]8;@S(47?>IIa2/<\=Rg>^<.SIdO+Z46WA<=[J9K;P>\)?C:bO8+5=M
\dEa,QPP)A@BL_f3(g]UZTb(B2\2Ug20GV:5,#a1F0ZMDF)XPg(46EQfN>d[\&MB
\>=UY;8bQQQ0a+:ULY/fOQ?35R,dX?a.Dfe<Ab5&X7D]f7gCRB/,<1[c^<]K^KaE
g8gK)#fK@fC1J@#SIJALcN(]bV#eFH8DbGP\+Z5_]K]7_:cO,4^DVScU:_^@WES8
P;dO#_R@@P,_((9]&RYO:0KLQ;[_Y-Ga4?7PJ.<\<CbL767fGN;b#XG]][;,R[\,
=KcC-:ZCdIGf.#\M<AgB3=502(JHdOP&@^bdQ_-LA?cgZ2b]:?J+?a96F47:COR7
<\cK>(.R>g06HQWW.TVg(4]f44)dUO3R)bW6ea:2XFGN/OQ.D#G0e]51+0CTJJ+8
XLg<8b[\YV,KQQg^(()X\-FIeFZaL;b3A^_M,@g;RR=S24f_(f;SFF>:RDWDLf:@
6eYM-Z>DHX#QbMS6TWd1#@K#JR[WD(]S9:D4.dQUP2^U^gA_A?d^.f2&5UH/<,:O
J<DT@\JZJA(2)Q4,X6\(DJ3O)^8Zfc-Z;@;#+9Z@>7:T;]ScN>N7\KV^PaeV\50N
OA)YCV6eVFR#AMaf9(\R^=XK_b_Z2f@ROaOO1MG]S<4[,K,Yg3NA,#fOdD@+d//\
M^U@EW<RW&M=T?;S5X8/DX2>1>/:A)#EKF--#ZAJSR2]486J;B=J\YHg8e,ZH8<.
_R#=3>0?I7=_N29I5&:P1;#R12dDMVKRTdL3+TB=QOdNJD;\[\9f>DZec.F>1\\R
)S)51YKeZ@JORdY<AQdLD[>MVMZ1S\>-I<6f?T;#A<1A+TM=H5a[B:Y=\K_LHEFX
<4^=[Z8FY4JZV5bKc]/&IL&360)FU?d15F21RXB;FDH6=3KU^((gE;cX..VC:U;\
U\+ccC(^JKCI5B6EE-7@YMMAI&4L\;-:d8<[52g1&+KaQ,a.cOPaN=BFLcb[Ba<#
[1MQF3(HWX@0EUA8/?Z3[+SgT2X<;&_(0._5fT3@45L0[f1?Eg6)NSd5_-eX8Y.^
dbWW9bWFa2VA:E.H+FWfN<Q(bG0KDB-8c2Nb#c=2B>8<^T:e+OV3Xce-<eN9;,L;
E=J-ZPJU]RK\WJ^aY?=>8UYZ,,F_e&\4a^J:HEULS]@&+O.B83M-C?UVA.Z;+LOX
U7B^6GNKCL,eY,O>.bW:-==(#1UU8]S3NNEA#_U5bQ3g>F,.0XP#[Q7WB1+F7?gB
Pa656_M<(c21:a+N5KKE+]ZVJab<BTb66O2J2,<9UbG)cON)60eRD8:>U-0UL&@Y
4&b>.U3VBe[8B&RVA#ULX32>A8?;FJ--51OC?];K1((SYELP)=T8=-dI\SN6GCfH
COee2f(QRLORDYe8R?P[:EJ71HOG4.&#/1(>=]:1JZ=F0[726NR;\b6fe=CO_M+d
ddL9:<Q4@-/0AaA<Ve<3R[9_?B]SE0V5[+g_H7E]VdQEAGae#J5^W/8c-LcM/?T2
+K?_C+bb>IRV/KfHJ,\)1VE4/DVT6L<J&b&1CW.::W7DNcO-0?Hfb,CKZ/.;9S_d
CPg;A3a:,?MASQS0QFQE3:2XFD.5S&<:=1VQ?>JD2(K:E@IKH?_DO.>8+YY+JL]g
);=TH(-]I8TL5d^\N6T2K^\8;.b#_&gS,Z\+a0L)bg6E@b4FQ0Pg);I3-KR_T?Fe
1C;<Se13g)QM0.124UE<>ePL3B6BS4[77FI9H_4M+?C]N3eQg/&?IO/75_\.]]CP
=22\=9Ra8F>35R51]Ld?Z/6KY)c2&;Wf5-IU9++84AW(=WMc]#].Cf8,.+eGP@a.
H\,L4<?MGc0IYOac+U:faI^DK?-;9-_fd\&P4,aaDEdWb@R-CI>HY^UPZY,WY3b@
),UUfOa)C9M0\-f_18NZ/SK)fT#0;Zd<8986B.O?@=;S.L[D(9A#.eFI6WN>R(<P
FJ_ZK9V5gM2#Za\(B6bdC#a.JX<XOfNeN<NQ@MR;V/8d_8HRRg7_a1X@9eM/].(g
?R#Oa6N/_b?4Y(1FC2Q<O[=&/@-ID+?dZ/aB1c1MD@gAEAFBNHV,^1OQQa1UM#1+
MHKJJgg2??bHMMD:[?X\IMDRH/_fc?JNJ?S[CcBY@#<Z@^Uge>-#f]:DHbf5L,_9
K:g5)NF03,\<KVY1RXNW7^&,UN)XN@7D^ZB9?YXAQ[]=Z_POVCEc>\G(8)EbZ(4J
ULSHT#85#(WY3Ke1<X=cW?28H@KM35@VMO9)A[Z@DGb30BKU#5K@X6,UMZ3)-(C5
<X#3Dg;S=JNFQ]Qgg8G0PTG:W]UM\c@X@aa0SC0BI_)1W5K9_J/4[@ZFP<^Rb8g2
ZbQK=9;;gH.BAES(,M/3O]O^P?KRI+(KDU838]&/CCQ2E/5g0\IGS+UI?8<@R;@9
Wd98E_H_1W^bg:J7eGW>:13,5>Lf-#e>X(Vcc=9-:)T[.CeF^=(>@UbIcWR[aM.G
##7&MJI/Q<[C_X7C1RNLCZ3ZHFc_H(gGMg]3#F__]f]P4NRbE-]V]](81DV:)8Pf
.NReDUZ<N#R<CI<^SH+EfKJ&XM:3eK_IfC_Zg#UeE4U/8\.T-T=bJa.TBaK[cAGS
PM[]D1+=]IcIe6->4^R:3G0g#+V28^L9O&c\W/=I3X]5a2Qg;gF/45f]][583)Ig
>;I&d.\MSMMO_.\Ebcb&O#2W7QJ;]MVdNRN2[]/7_M/<^>J?9f_e>S@9O&CKg1KR
[F@ABNYP]=Jg_,a5[9b_?R:[ANV,K(^aS[XTSb(C#AQDNKIH1d#;SDA,Ue[HIMWR
X[4+1MK2;=&61Q)S#(Wg)UW0bSO4KWEa;G7K&bFaGW0Z,U;I3G<HQ7G.ROA+I+&_
eGQ4SG-M#fdY6005[f/I((DLE?gUFHW:BQBgS.@I0gYPY_g3?J]aRPD1C_2PA[dM
cM?..02a,693SM9L9;_?)eSL7d(Sg0NK0b+c;OEAPBR5AGPE05N[V1=D4@[M.MVV
HCLg0)A,X(O&IVfY>[4DTdY8bJW(0)d[K=#S=588Y_9>,c0Y+#5O[V3G\2aY4aG+
(GE4W2(^[e(\I0&2F.d2@3?3.HePYH+/0.+4:XdZg(=)7A^4M_a(3Y<P9e0UVBPY
HcGQ(D360)DYTO[DBPGNDZHCLGNd)Y)S7[d6_fQ8/1\=agE#25Ud#>])I\BAIW5X
<&UV3F>7Zc/T_90KF](W9K)gbK_ID/02,cK;>34cf+CUY3L1W:_A,G3^]EFcC7^9
K)/Q8<_A;_RH#PMMTPe[^J,F_&;1fJF3CAOHfJ>02):;dG.eVg5.Mdc.)M@3)#ZS
<XU.Ef\<;XJI[5Y\)J)MH)+b(IHNeAeOG#b)6:MBKA)K3R7)D,+G0d>MQ1IX8BM;
He2RNfOG1G]7P(3=8C3CIe=WGF._AQfScP9MSU_@MH(4^aHfa?ZX=QE7A1?C^?Z8
C,Wc]/c@eX+L\,QQ6[Y/I+&T3e\&=7YZ_S1G_=8.PFTVeER-^CPa\UD>OG?RfN\(
V1@g7V,,.4Q7GSeL+FOD).[JWU3RK6&bALYb\IM4:NcZ-18R8KV=83.]BB,:3>WA
ZLX#WOF&]CZ@Xd;]X.C>Z]E1XHR(T=3N&Wd^9(20AB&:=2&aG9,^&+6JHZFG,S@0
.d1?&YBgGB?b_ZVTKEY^4_E:),X#28ECYNHL8c66aE&IV9,]E<F10_=A_>8Vf?G1
eY]=gb+&QE3L)2Kf[._HGY4\HW@gf>\fRg>DF9Mg/Zgfac35-JeX0JG]6;1J-8,O
8B4.a_d2I1/U-]?RJX#c>bDR.O;N+R4Y?(\(FOP0FW@FSReZg=/<G7ab(KV6IfNH
5KHJQA@PTV]7b)3>RJb.,Xgdf47&aDFMDQS^R)fK3,^#KW&Q0OKJgUe@Zb.JU/B9
(SHM3)HD06S--Ed.\@a;WQ=@^T<C05L>RLIHUJO.YUKED_a=QE\U00adIa#GUH:G
-H+,QOI(P>HYY^N3?dP#+VBQ9V7NJ-J6]3SUPQ_]>Vb,G-83+KR=LfH>F?R(JVQb
5,A@X1(Q61YY5Hg@64T>/:#0eQ.]?L#Y)Id-[?=#[Y#GMJG>F)73)Qa@3.[?W1;G
[4,OY?.7LcNXL7cV;/R.RCO[c,J?Pc2<-UgK1Jd;TJ_+)R^CVc&5D2-.92=cY,W^
dfD(WcEb6f&/-65\S)MD?Z,[@f&BL,^DJ\Rf-\U252S4bP^b[K@4G<03<2TWcZYd
V7GM2_3XSF_a=P^UO;7K)0TQC7D@U,OOC=]60WSYDTP#+UQ>&E5&C?R5cC&>XSIR
AgdA<g#M7aNd5SULG:D/W)W69]/^@d^)-HDFP+gJI=>-B]ZF9dEU?G:CU.@c[3La
EEa+T>3HVFPWYU?;?E8U3-B?\+#fVCX]NNY:V\6Rb>[U;_8+#K&ILcRg1b1.)/G#
:/1cCP9O5A+<2;>=e</-K2C.32cBYHBeG&;fgPaDJ<e=B0I,LLe3c?I2b1][8^7>
VZcEN9U>1+B6.f/X^..4[BNALY^O;M?dS)4.G/dLJd\@b,EP41f7A.^BKQX7ZQ\f
2@bJ.D8&A8-]dXS9aLT<Y1Qb2IU,@a?H.MD>0UabAd^_Y4W6YH1(WP^,b>3f6[R5
DB_0CcL(\E_.-\<;/6#3G[,)K8XPdC.I@,-@NN-86(_+b=Z96(?L0KW0FST@</cM
.c+:)0PH94?O#&eR6e]B&/+&];I@O.[)d+/4aOXSV_Z[078cDP)+:]dSE@Z[\VLS
EOEE_SXb;Q+BMa)5C<KG1dP@/OY.WKd1Z.dc?0:6Q+N8gB(JOAf+70G=/:[ZcH?K
fQ(f<Ke8?R>b1NE=&e:G/EIM^F^&_Yc<Ee[g+6#R8TTKF9gS(fVNEZA-VKg4++D1
c-.PA&[>OI)WUXFD/3C1T>KBd]XU?+9dNI71KJH7]cC_4dPS;Y(90)M0O4V[[-75
:WH?Wa8#L#=a0ZE9A=AZN>PcG\C7\&]VUB>YWX@aI(V44QM+.5(M;[D0g#b1>Bd.
.,Qd+;G.O3#7\QcU#Ve;UA:b&(Yb.d=If)aHUgTWDcYAH_JSIDL\P+-:WIbKE8.Y
0Z@b?N90+4?>;DI:aB/5P.#+2EGG5]6SGK7[;C@GF2]5_RUS:I0,^G,K4_aUV@^6
/@.c/7>>7PA<<Z5:MSXW37[V.<;@,(/+54G(\,E@=J,G[,W1V33=2b3)@G=dd>0U
Q-:7JTV;f<CZWdRObaMgROP?-SM)_I_=AY&,KH,b==;4Y.GN,GgdO_7;cHe]cBgW
#(Y+]f<2X2TBVg8d0)<7215AZ^<^^^IcSf#/+Wb/aYLe1CMc\&PXV&N538;;.^9b
Se#NFLc]@4IW@149\EJEFdb2XR\E=CNVN^f6:6Y7S1R.5R.8_8ea[(bc.<eaVOQI
C?M[WK:U#_SHA;V7HA:)[+K<8>I^O-0[XE#W,N:Q&[14CQeJPB^B1OAEQd7:6K=c
1_1KST#EbW8W0I6D9TAOc>L:RK3XVFDU#fYK\e^H8[ZWT2@YHXAN+^13L5Y,<SXf
&=N\&D>,#3]OET(YfDa+G74\YD9[TIM67<M,XYON@CVWV4eE(>abUIW0bAf2))&M
=JWGO<EH..WAIPXJ]<dKf#7^,=>X5A&,Ed@TcWXBB8ZVPRSfY6V@13^J\N-Q\BH/
ARP/XQeB1V296NLcf1=0^f<O]UZM,XX\@eO^8DSV8R^A;#&N<cUZ64a[#?K:AUW_
Z5D/;D<OA,^d#^>LV2[Z+HNIX,W.C,9G:19[Z9aHLSCP9+34bO]_?C>@+4=Y(C:&
:C+;,P05\NK4Z14eW_9c;#dX]/^HH.&D&._48QLOF8UdcW.0>K^&6T76]JQK=DaT
(PY3@ab(3Hf+O._4U;7S^<(&@Z&9\;b,.?CPdZK<:WF+FJLO)_#CEP3dH>3OZNUY
[>;Y1LV_g#1V:e_S/L,^0JV3:FV3^Rgg:9Pf&)^b;<7(BaIX)O:#8^CE/)AO3A:#
B:Q6gZL5c(9QFH(K\.95Fd2_.FH_WV5&SD]g0C.<eUWZWHRb]>6CO&]U:RH;TfV[
;AHQI@5b/>/Y,EDE#&fc[3/&K?\\30KB1C1?I;7Q.H+2K?a?\7B7E_P&eQ^W>c<Y
,f#,Z7X_6_2b,D4K@3UV>85fI\T<0WW+4/&0EQ1OBY,J:N>Q&8T?<[>b6L#V@bK:
>ASRB==5OfcB#OH8;G8:dK;/8YOQ+TdQ&>2<<Q3\>F9Kg.8)2KKc@#gN-LIEW#X2
[3IYaeAU,TZMKXB?HdcTMe,CVR,?DL1Q_/PJB4f5Eg\.?+O+_C/[AQ,4S)?FK,gQ
8-LYOU8ZL,-d+F&6(#@&GMP8^V],WDQQSg^KQFa7ZP9D>_S4?WLG^A^80(PYfAE;
Q2L3#aAA&E7?P([)e</9dTL&:XJ(Y.CfX3CbMI(IGLaecLTf9#JQ-DNYJQ8A6c7X
<ZV9X,_Yc\b>D2SD-SDbCX[1F>bEV94YM5E+><V[@G6A5@_:e[H,cIf4F;3W[C9/
I6FWId9I>OMO8;GNQA-@1T@4(9]aTEg?;a6gL\[7bAQa:@0/5\<:=bf3>W\[dE_^
CTP?Xde<.V\2S321ADE)##8Gd-C4)[5f_E6KU6a7?:.=TD8_2#QN[[@LGg_Pe:Zd
ZPBe1),B=f(bJ.4.84d;:.=Q3G-@3-X(2Hcd,H[;][V.cXbMOH/cD_>CbdJNR\B[
9+NS/<94a=Z3F9UBP>01aBN1XJLe-c@YU+6WMUR+^JI<GXQ\UXe(10PUVL#83e(1
4^5#gJ]OJ<4#H-ZPZ0A.L?71]dVA\(f+[6-0e(KLJ^A,(T()D<-3HbMZ#:+WM03W
,,=4fLIJP/N<51f:7<IUEb#Z1IXVWO-;@eK^XK1-^+^^cJOVC:AOX4M?(EKJEV^f
N3aUQ+(RaV-#D/Q=6&M:HJ>P@;JU.J=LTM(BKSg;@IDI9eA#_C1[-7N6@@_-?_[b
bPA<0Z0)8_M.FM-_^U2]2TQQ,?2RU>19W]6?H91U]dBO07J_\&XE]<:+O/(b8E^U
,REOD&-X;U(]JMcUF4(W6\7E[M;LfXB7Hd-Y+-=eVd9)f=KA6bd&-F&JU\(VL19;
J50#;0eR#DL[[?TV0SC_>A4F(^PJb,S:K6Q+(=FE3S/Dd,BZC].9-aXH=g[#g6c]
A<HfQKf(F80?;9g1?IK+</\Z4Q6Q0KB[8)P-D;EWf1YU58]cS3]F1N8Z(.J\:/[R
]N:[.=PN(51F&G:2AR<+?@H>6NcENU:B[0@5T:Q:W4Z^PXV657_-e30DK8=<#c=-
L?9C1I+a-fHB=BSD.c]ALA@CB\2/)UdfFg#FKFG)g#NUAPf_3N[(R^aJZ@^6:8-N
\\/6b:G:^g7#-?&-9YJd5H+VLVdA?QJK=Q<MP&5XNJYC,@\E461H9B&8L)=H)7H.
f:#HYE3Q)T9e@HA53O0N++O2H;a8;#5TI]]bV<7]>E5fgCBQ74-_3&]F]M]cC9^0
ed8^eb7-B/Jg^[V;^[6O.KLgUKX_-L/@MA7^5CBVEU5-42/+E-efZcC^/H02Z@gM
@_.eFeJK/VV9M-,CgOB?6B+1?e?^6QRJdL--f)Y\I9,08YK]JT_(1S_@d@BLVJ[,
c,(2IMa,3XQ1aO&,36H;X>N81Y1O_GZNg(V-gZG3))gb9ee929#K_^<)WC&8OfSD
(XN)L5B[EHH.>bL<6S]gD]W/QL6ZgG8ab_TH-+MQDgG/SQE6CHV)V<;\@07^f_KS
W0OfTI9<.9BSQe5800K5aNLgYQL8?eYG@\<41C,)17e(+4IY?Ib8>faJ6b-9=OSC
3S,0.VSYSFRE[>P&BYMHK#fWY<S//1NS&\A1c\FAU3[9>17&BJB:fLVM8Xe3HZ1K
TN:f^ZS4g7#89Y4DJR;E3eCc/LZ31Rg;/]_=49]LIJ-9eB[b>N&LKf>6NYgI/6c,
-g)ee\XUQK>1-a#f,_aI3.ZL];CgM5eDK=O=8P4C,<.\S1/1J/7CTVD4)K&X_AUf
1/SBEP-AZ&3R+ZC9MJfF5\[a\,Vb2BRg17A4K=c@d>MU_>N8Z3JcC:(F14\5YNHO
<.aP@B_egd:Q5#TR^74[)-Kf#:a@OVU>gf5C<A3H&7JK-]#d+TRcN,d1Lc6/DD57
Db4TD4?0RDH7Va@3K;2YQYF:MS(XU[cC-6-B-g[\)V+(&2af#(^^C8F5.O)3.T5#
Y]2NCfV1VY3#9QA^2H88(\02E@<bH(@Ea658D49B9N?7BLS+3#b19?+9M\Pc/.@U
NCPE.d&N@C],+J3(g\>Q7B>BQ.[]3.V27/D408[M#20[eISN@/C.JO<\109,O/I)
@a<BM7/78d9DcB&&/>AZD-fRADV@Hc8E0^dA]Aa;@X_J.SM(Ve@e-]<@-Z3&D]HH
.1GG_>)G1EX^E)K4U:W0gQ+P<KDC(eR10XV,DePaebg^d6\:[0]M80,g_Z3D^+\L
a\[NR-.efPRQ2I6BC44M>)C<4(:Z=0.K&]:TaUB90&F(3..]&^0)(V9G:W1./b<7
>H(g<g^495C[eaC643GYEJYJ8=dKaG[HAa7L_T7Bd..7^PMLI#/P#;I6\VT_X5^F
1[6S>5CJ<4994fROE)7_;MZD>)##XO60Q>J#3O+U2ZL,_VYWXf?2JA/g1Y@RSRgH
4_?HDQCb[1)\X<YJ,4]FFHX;>G@da,?=6A37O#K#K:TC)TE2>-F1CO;B<?b7fXg.
b0@V8FdVS0^QO@BO;eP;@G0]aDVJVQ3-7LV56Qe6.W/gMV42DX<^@O^@^<&O]H0C
DPYa5=ZP@O>A&IGE01SbbAX>Tg.1eg(-eCKDb.8bT<ged;/CYcJ])U5-2N;77UF+
>7XWPI6D]5YYQ2SN9PYa3<B<+M^0:XcR)dY#aF.c???e8+e07?U@(0C(^Le?abP6
=CJgf@5D/2dHQ:)J]#K6e,aPNTH3NH+_/\H)])I-\HR.Q4;CKTb+P7[aPVBI,6?/
&:f2D=8=,Xc,Sa?DUb:V1^&<ZeQVM1W3BHV_PeTKVIVLIA:Ja/2+6ZA65fNUG7]R
6RbOWb54[LDMW4Ga\K>cT)&4GG29(<;;]_G_b]2?D.C421\9UB0CT+?e7a>6fd2T
ZcBVFR;W56NZ>g&Z.;0T6L[J+ROO]+cVNHN8\^3&))QWD(GP9T4N73-[HR[Vc?2d
BUC&4SI(:0L[L7=/Af(E-=Ha?AB38E&)F(Z,;G\ITWO=M,<IBD+e2T/GLc<;S/d4
0T:Fe/^KV[B2N^D^]RT9Y2YC)6BWc@<K1QdbMVCbg+&A#X_ZBIPGO@FCA#[DS7[\
56+0GQGgb6W?<TE0aFZ#66cHNOD]IY;DEg.5:,=,9JLEgB@#fK7d1].5B3aG]PXf
a@(HB:9dQg5&5?3NMC7HIR1#-E/_SRZAJO&DJ94SAC._I<B9H/IfX&;[KdV^_7fJ
\P]eVF4Z5FKK4/Z^;/JPC-H-fY;Y#ZI3MeV2^^>PR>OPg0I&T2Nd^a]U+2#/7YH<
EaSA=E2YN@>;a;E6^S^.8IW4KYKHV=15D/X(E35;aSC]]/Q)Z3\9KBSO1H.[1G.Y
@P^9\Oa/3c>(^QM+0^PJ1R>/-O@1),0523Rg1JT_=_dAU;<A#c;\eET8X@]UUFF_
QA:#YS=10g25EO+VB=7TM;>NIS;Yc.(#?fYX3Z<]FVgGM99=cZ\[A@QgeB@(<_B5
(()39dG9<.J68UYbQZcb3LYU=F34:^R^36?EQ^Ga/I4M2O9K;_c[g.@#==CB7MCT
TRDV3_PO]-W>HEb2e?4FLX#:B#Z)ED:BNKL^fe)>A+H0b_-?>CXR6TZ-I[2)4P8S
X_?d,U.UD;?\.DT9-#JJO&S^c:[N7e8<N5M90IX+&=PgM0>g@cKN7aa&L>JRXf_Z
RICS6-B@OO8ag:JeCbCR8U;5Q2:X9Y;TKc-J6I=SSZQLVEWI,\/8fcL>C5Fc)(,V
86VeH6e.PAZQaTBaVP/Gb+=e1^&3G2Q_Ig2aNfIE6<MUQ)XPP+SBeR@0G_ICR0=D
F@LeXXZP1;(GV=TM-NX)gO<&NV:@[1a/[Y/#LFHNd^VO&2e,a4YBXVaeV+95A/9e
g20+g_TC?ZD+/\10_U?))_>O[5M)8#g36W<@6d_>=\/OH[e=+>2R]MgG>XWf2XSa
R=O@11[X]bTd(:0)4;XcEJGVAZ&I[8T&8E.P0:XG;5BQWF+e@aPJ\(ZY8OF0+;FO
O#A&@&PDBfP3e2Z(YJ\gLT54V0NR;cB_Y<2a<(ZJK#)\#>Q+#&#768fMg;W@PQ?E
<V]aI\_.H[.9&W+d;YYBED=;-&[62BbGO_c2D@bMK9bKCMeLFA]^#I]T\DgMTB7L
IBTUBA\D^H0fNTR1SZ^e\@/c+KO.UE?b_H3]1&@U3DA3JbQ;>&C_XDA)I(=Fa8P:
YT[B=K54IcEX3d9VL_)42VfDG\F22,09MGYUcHc:SEZ06#<2N;G3dd)g\,2E-X((
79;?HY7XI7=M\^X(;T#/P]4^SW48SA_K7OaOV+]N+&VKLH2ATP:>0O;BW1IM8Zb&
1<:2/C?#+:2Y&B]@7G]dB>f#,=<3JYALO6JN<g<@Db[J?Ta@:e;#AGc>(6fQDP>_
Z:P2/C;1^/B9-<4bV:3M92&fK98R+8@Q9Ba/M2[C-/_>+5<g-g)dc7gGOB-[,M60
_F>;NBHS?XXHfEBbde3GWg?M->TK,29c(?(1UYJ\NW_>UfYY@GEA4FSPc&LE8c0c
dERYe_9Re&:9/C/\F_P8>8.a8@TRSGS0-O[EP#Jc1Q^,cZHD.)0fY2?R2M:S(9#f
&&aaE[:71;#:>dERdOX2:/\e:GAZU9-KBQEAAbJg4&NV[Ud>XVA_11H\JQe?BS+c
Db[.8@L@&HQWG1Q84#&EL7AaL&PKL-0,J=Wf@VGB)60Z;9&\7[\fV6XeBZ4#>TZ9
]:2INP63YdL2276Z8d@P-F_c&N;1\MJJ9>cAZA(]PI7M(]+58GVHH/+bVC#HP@4+
Ig2g&KZ<OLa?JRNC<A1g_dNSX+MaM4UH4f#_IB9X86a=7gfOM3C]0Z,_--KNDgFQ
G(>N5L,4=bfYPT:TG,,[RB>Z3W@?;e<YaSH+Y-<e[F^28WQbSGVP(-60BYfCI7;H
GSdB7d]\)c=R&5,]VFT3bWaL,>SRBIOJI5KT,DXeV+VgB>Y\XXScAYZBcgBfGC,g
(cC4TfFX,KE)A+LV5ZXMb=2B@VeJgEBPbKUS@-AC2H.,XZ\?\[6A_AM05ba-<cA[
^(HBZ/?45B9@^5Ld&\3VU83.EaaO,-Q[25=0&bA\gf2V:a]<+N[2])a,8JIF[MEC
U4DLA9\FQ-K&dRT,R1(fFFX9G]GH?a9f,).RUVG4L4]b#>RM^NOLUO1F[+QHIKF3
:CT7J9BLVB<K3.QCd?[FQ46N(@;7P[/[TdH^]X@W4B?<dTI0,G_TAY3abVU(@-AU
]NT7Fb()#0&fP5X4?^Gg>]?/5(K7XMXE:ZBg@DUg.]D5.A[4WBW^T[eU[T9=aOD7
686K>IKcY2TW@-gZU8RH>UO#M9&@KM7631:TKe.T(Jf?S;PbPAR.^)NGQ-5gfFPW
3)M3B^\@/R53NVF+#<1\]LK?e9)^]NFa_&BFb]dUc[GaOS#HAA>EKCJM#M[ebY61
=Z.Q1UF9dG)F.GQe.T^=E>OCVbK<>Xaf^[&@K+(L1f#I[N_Y@ADb=9ccTE)8Y>@9
F[V+b[::g]Y)]I<g(f;3DKHGb]OcNc7),7,4gD#@YDG/)BB1OI/&0Y=SCFU^2?aV
a,[#O,1;D.+,]LUN=L2C@NCVAXLR^@\3EGc.)B0E/D6V)fT@:C1g-5:S4JQ3#&-4
8V9/4IW^XU#2AGB#@G47<045D_OF(484Z?#aX-6IC.T?QNSR1-=b-J,1GY1S?&[H
A=3<^C;LS-UIP^(A].c&D\43UEdYQ@Q21PZ#++VbW#P9RgJXQ]#7#PfOVXZLd0&7
JO6V\/A.P7W60(#BSIG#^a1>;>JA6-J(KacTB2,_VGL4f#V&4eZa@NU_3:-R6H7f
?@a&:F)REM>IK.gUJ-G)78g@H4UN,)8Q6XZ)&9ZR-V9(5>>7f4g/c=b<WHfI;E8^
XS.EbNfgDB_#:I+F1-&SG(2Z&NC^aLYDFBS5;9N3/2V;X7a=N2-YMGVY1\&cHER&
X0GUSK21K.fC7;#NRJ@eH2>:<>fDL.8^E7L7N^\/YQPB#5\B.CP]Ea8e;X7VYEQf
T?BM-;6VPg6=9;O^WS\=4(2Y^16XE55+WBY((=;<_&DcJ#a0AFG^)c(Q^]#1&W1G
7-G#&O&GXD6)##AAN5(_4DgH8fXdP4]SMEN58\I]U15Qe51.C6VE_>WfY;,I[C6&
B2120TG@+0OB#bF:C>Ae[VT0;0C]DD41)<96P).J+-T>U@P;8.6Q_13PGA]TRZEU
?a&H=WO1fJH;.G3BefcJ]Ig.J_]L=H0OLG^]_C@Eg+CfPcAeE.9VG&1_NF/eBIEY
\g,5fO[TYa-K?P3:&OBQZT;1B3c32Ea\P\,0>KG=e5E?[V5@Jc2/ac?[>2aOa_L=
,AF4WTJ8Z??55bCZGXe)8>#E1?a:(W.4[bFLT^Z#IWYKdD;QD<\d?5_Uf^-WKU2N
6,(M#LKNa?=<+O[M>6[.P\T1<8-PO2_E1X\X;G6a5J8_L7Ef+W&620IW(H&YZb.c
aCcOB&?04VAP./VePG3VY^&/VE0ER]YJM4E+([6XZ:,YbV/de?fbRB[<S&EBa^E(
cIV_#VDS47[+-^ZH=:#0&T4(54.6>4,DYLYZ8CUb;Ac&_WUC7_@[GbA@XLK]8W8[
GdL,/EB6f;)T_3.O_^aKLI&+IOeP05E/7\9DW]5YbDPebR<B<SISgOZ5N1WF@fbG
P2&A0)+A/X3=_d?E:cNJBOUX(^Rg;UI:KK-M,(DB>5IDU99V2RX2#?;LbX?-1F)0
YYVCcQgXc[7HNUTYO57:0>A42=:?RG0JNPc1)+<D-7+21Q>Ya?7YH+3ag\5RM6-N
1Z7;\.G2LHA@#2)4aU;M&-O=IEP;/Jf)A#L1?A70TY&_235Z@\9M\W5^:2Zd/8-P
YG1]#R:^R1G?X=?L4Gc,e82)CcH&OfR[gJ@W7QC+Nad9e_J)3#Qb92cP+OI.<L4H
c\f808QT3Z1E=LOPJV4UUE=fF:gV#O4,QAf[7HOf-QFcG[EH(XK3(8;^QWM]d2CH
@\bCJ4b\g.KJ6IR2g>E-,+<Nee:?S^7bB5VHLK5)&O;2.2HJC/7(W:g6<M2@A1aL
Q/:TW1?14eL2WN7/bIc.&3ADUDNbIKP^Q)NX3MTU/+W;:>-6[BANUI8c194?7HDg
L9L;6OXe9(6f&72U_?gN9Q,ND\6c)>N8>#6F-IUJ71F9b,^S&6<GUdfIX33L<.R6
[aWL<,g&X0(R),e<&b@]BJG,,]fdOAD5E87_43AZ7Y?VRI1=[X7gK2KZR2b,SR0@
Nc-P#])@@HdWZ)<]C17_1bT9K9B)584d8R5O<dK.P)2&O@F5E1;5[:-\8DD,,Re_
1PA.Cb^XJgdPXD<?&_KI2RP2e-Y;<Z]9_2-9>&6+86TQ+D1==eJOYKG5dd9L[d0e
=ZEd64&[.gf8#&0?SYAd89R_ET8,7+0:)E.def<B&BDH-><AcRC&7;E.G+.)SaL6
K+AUAV?C7L92CKBD^+VIU[4=M-]HPD0;\adX4G;eAL3f5ZE@[BaH@D<6<62UF#QJ
0TbRK:P[b9G8#:8N+;7>LFf@Y,G0Zg<Ge72S9:?A9+bM?b7#/+EI6c3WUPfTFSbM
f:Ea(-6DXV.eb,3W3&Z\G3eV4FBDUQYZU&1fZZSb,YX]0BQ(8J]AU2BFa-2M1]O.
R@2T&B7PYT_AM6d_N(#=KC#JR#eOX0cA4VaX.+W65cTSJND,6\?T/;7N0\ZRL0.b
BJQ0V3#4DI4]=/?:^[+J7/J#I.P)J2>6eY6AFW8)PJU-8.DY=IY8Ua]ICTN<:C=4
Fa?3N,XM0,g7H2f3SZGI9bWZ[F&P.+WeePF,CAKE2/2NCae?&+.,VN<]\f5gFP3]
G89fBH\YD:@F93V)1Z@Q2XUcWU6e:=2=IAf+X,EIH&dIeC]FH<@VNW6a[FVM<+O(
6FL4-U3,9<M/[54_(#6;.H4C\OdUbR7N.&KLdX)49(IC2adG;PJ;1N6Y.d5<fP-d
=<V,ebZ]ePT)9N\f59<#/g=TSB36>R+UE;S/1,+ddK2.U<W>N9aQ/^\_R8<dLE?O
+f]Z9_\\D=T>c]\B2V&ZEOF]8TXSfgP@5^4#7G-g[/5P?.JCKVWOF\PNT>FU=T75
LJ)?31_O/@([I[5+d@.RGQXLg6;YM\6HAENS4J/8#09f,76GIN-A6?S.F7<00?</
4C]2Q=UGGMFT?F]O9KfMcF4O@=&9Oe4e9a;FJfc[7cg:H8?)>4F,ZD\7J,G/21+e
83<\LB?#F\We^^?>^+-8PE5S,T=8ede80g]BR6\=H]BJ;MCgEZd:LeP8TVbCXL4Y
a^?VKUTL:A-X9DQb#LE^ZgXVYO5)O2/]2Z-CK18>Q><U7)e&dCad82S).P94A=g6
TZb4TU-gFM3Ce-b,5M6V+-F&5]Z-WY)dd_=X(H=b:,6a#R?:E8&b/HBT8]K^A/8.
CV3XCC-eX3K@UM9@DG-(UE;#1dG[aF(=O?F)>6I2Z@=BA+gCUS0RO8+Ug4<_&H8D
6MLY/)1ZD;^;cEZ;XPP-L3I]@IG,TX8003P87PLX-d.fU[FA-1]1caH^]R6-G;W/
<5>VGX+PQ_,?eFF4a:A5PBBH)YBJ&AgKUT7WN]1]BRQ;IZM-.J,c#^(e==P<VO-<
I5I--A5b7QN\;NH>d,;-^X3=-I_1RbSJ1g_S9-1[0A=0Y?G0;[9#&/J[5J)A_g/O
\\e>=_g16a]:H=8K3cbAX3aK_./@V?[YB#P(P[^Ue:5F2047.6H7QcNfNFb8Lc_4
.TBb7f,)=IZ(^SHNX,dN;6-7cFbHEb+YMX/ST4Eg<:&MebZ=<YaQ>2NPXAECH@SE
/Ec#cZHe,)(?]1M+31U&]R@+YU#B\dQP#I>c0G_CNKd5E/<2G(HK\?1K8]ZD]cJe
\Q+^@BKaTe7SU6:0[MQDXEA()&a&c7@gNZ9e(Ee=CgMAaf,W@X(2)(G-G46U?T].
cRN45EB_.G7Z@B4=RGI)-B<X-P8/,)O^[Yb[d2OUPI([4YDVgL:eS)g62D^9daE6
+R?C+BCNC3BP7V_#D^e?35=eN<7I5XVH3?3M5[F<-gC)+,B0J1d7Aa@Df8SD8<TY
#)(cUPG;ARe#=\OQ<HdO[2?9H6O0e:-H(;\\0;C(<,-ANO6W6d/@1f#BeGdCTE1T
18;EfS&bFF]47?Fg@^MDf:&CH?9S@BF3LA(XV[JF3)H1(JSOec]b15SQ2CBeabMM
;PF#U,.01_eL4W?1d;4S8SZJ4FO@=44>88E7c(GRbXDV8CB1/E9/1La2c[1C2R]<
A9N&b.0U-J0/3.,]&a)g^?(BJVS[]\7HL?>8AX)RdW#9/^L)IgQg^S=ZXEWZ,Z^b
C2FPcE0Ce\,B^e^2E8=B]JY1?S?TH^=5X_1&@c5IIWP9d;6X\D,]A<&[K/-9]f^d
<_ZeP/3>K\FH>CU]GdB>P1a^;L<I_ZPdICDd[2(b+&T[RFD;cK0N@[999V#F1c?7
e.6f?F8.MT=f857@A6c-BL/VTUJNN>P:c4.b\\WAD=5b+SFLTVb@<8C&b^0)bcA-
?,]C9aD(I5ORFd\]:NIH9K)HDLf^BI];Q;,4V)CGF=6dTfN.]6#0E:bc[;Q>W4I[
5J2\0UK_eA[4EG80>F8]HKa)-&e-V>#KN&44/]M;L2/>/0J._:Q>#GcE7=CPeR(7
5QOf>D:4gQS4fTI+.&8KGNEH3[HWQT+9G76>3Y:21_+4a5cKN]-;^0.>F>0G/TAZ
K/)UNdeBSS-Zaa2cRSbH#SceVNX&8QP,d/5;PURdTJBS6_bU.Q<A8ZWV1f@gUIC[
;B3L8L-&\LQ6a5<AOA13/4Gec3&dJLL8&O,cP=5R/3=B^O7dfIG,e3/Q87&3[&H.
Cg^EREIJ?UQ-.V[W+G^9BQ@DEe/V/X^><M96-)CZf1GG[>Y_1W&e:V90H^?_+N(S
[SLE8J\R<(2\\,))F?ffQ5OFKQ;NXI5EH2,6c_4NaTX-Z&U\PST>c8U&2MLYXH#F
d-M=,Z@,ER&aR.<BK]P.FPDV(X:Q5EUG56#)45gTNZW106Z[aKM4IK9OePY?W0]G
8H\H:3/eCRFDbSA7++U6]]^-CKD8@(]d[@O?1c5+UQf#d+T5Ff>L]eK:c9ZB((#5
-LdC]QKbUU4]BIDU5e2];/-0Y<M9_J;G:[_/TESRLKcBZ2QP.Cga8UHNFDaZ]W:g
:YNLJ58.X;f,Pf(6HOBg>4KO8\7\IFX@T<Me/1d(;FW7eGKS^6J5MC8S;TKV<Va&
>NG;+H4E\D@d1#c.H/fXO<@ONRT_[V6?@/<<N9N?8KAEC5RCcN0R.DN&)G/S@=KN
BPG:Cg\CHTcE+RS38(/B4]Q1A6X(/X>D_g\UJ&f&T#WQbe&<5651\1^/REEPWIM&
3f99P@7X,MQXI[KLOTb3?I=\=2(4]M+H@7L)F59PUZ+_a#=(bR=<[Ye-^faEd;8X
JZ<UQU\V0N,&L7LA<)1]N[_:6G@d1?A:Z[]4&F/8^]A:#F&=UZLab,.aa+1Y(HYb
-FDggCSYd4I,XC2]bDUI3M<BBa1YG12]\1>C6:#HSG5>TSD,>;5e98f4RNTaK2I.
c:_@4c-N8c4C_5Q:\Hc:VXcdQ@=@:X3OQbgQ@(E7\FFH6V2H=#a:7;23HLPCF&8E
efVHDLP-CQ8Z4_?0XBVL<d+@PF4]aS\cP<-^?>\<Q[1.f1Z#0W]77OK,X[P&_GfC
M)U6B3WQ99Le9b(YJH#8b]4D>AEH>/dCDO&AL.dTJ9?:a5CF>O)YDWD;A:>?^:UQ
5JV@c<8QKa-D[A&\3\D>C2F0)]NSZN8&+Sf=4IL_(V-ZE?)A+HbYbd89:#BQgW,^
ZH=>ggVN]V#-f0VF&^_Xgba12F6OfVC^G7W3QS=ZHFg5..(EFBAb&^0EdK@3HCG]
YVGD_,;_C()L70K;XH-#6GT0B=[LPP;QLTZ(VXY3D#([BWfK##d;\4E>P2=6CW6D
>2^:M:<:T5=:,Y59Sf>Cd5;KgR0K2_;,8<U1]IV].FD_G?[P0>,S0ZW2107/gETF
Bf1gV&+<?4^SC-BQM2E,9b,E9:NT^7[L-)eA2-I5Ye.:cPPIG?3KbE[P].g\^N6F
Cec1.NU-4FXKPJR-6@dfUd._7FRg]gg@[Z?d?]BR05#3.PO2E)3Cb6+-[YHeJFbC
E7c0<LF2a1B=VId0VUUQgK7WMG,/[&;OPLd?AJ_<V&1.EfKT>?CW>WOCb&.HgaDR
+Y;?TTT3&Q(#f\<;GEaQ,R2=+fKG7g):Z6M[aCf;HFPMaCY&M6Q4.IcOXV,](QZ3
B.OCB)1(ef-[/?]6fY4a:;,Q7-R@O=LZXUQ1H,L?V-&bC]b=U(.S=UX-=EL3@XA3
afK_Z60(,_PGRA00+Y-SD(ISN@[<gRI[ON?#DEBZaLWY@L4Z/aJGC7_3K<-].6/_
-(LDS&,g@FN<X&&[SD],:c?cAE@3fARIOg(Mf[0Ta\NQa)+G\\M(S4:,KZ\ZU);;
/=5VI00&JB9==F^/.GI=QbDYL->W6PX]e\e0AA15YF^f8bF#V>-M+;eU3DR7K;1G
0;97IcN3+[?<</IRaP@(U1+a\L2SHcI(G?HRDgaKHOf#\H#=<&^2].V];9,229DN
KZgNV(I^H.PI;M208SWVaDg_04a)bRT1>&W5LB))C7\]6FIc9^BCPVDb,[.Mf0IA
g:5c(f4^19>1E7TDgDTDU;C:F4>4f^MUQWY9MF^\gb453c0_Q0==VCZ>+AF:)@X3
8+<b131eTP[BVZ9Q0R&3&WPKCLN.+-(3:;D55_3H=+TG-]_2bf.-,2O9K\T&UA1N
;A).KG:-cS#JKIAQY2A11\(Z_KXH6gIZH^->N#BZM(?3Wb-U\8/IS#gJCYMf:_-)
))^RCdDKdO-.5d<Y3?Q2H=FV7ITM/4beI_=Q.[6&)79W>AN12N>?bJEV3]R_)Y)R
Q2X/Yb+Q&0;]gO\,RSV#Y]Af5E3X1B6YL-L:UVCc8M;8[9;L>85H6O-=8,Y7&@XD
O<.g,XQ@O#T].C5VGAg)D^a(G/e/0/H/3U]Zd5UQ.;X2c29[9(2Y=1N>)=Q6WS^>
9Ug;I?IDM<1O<W8F/7+Y6Qa]b\Q?F3Y0(XDegYS@E0HDJcXZ(]BSB;caUQRH(X0I
&:]FA+8ZD8b0OKW;PV,^LXC((UQQ-?/faaKQ+PE+51:A4(^QH;>.?<.g4OSV2/9F
HO;S:Y9H,K60?4Z4K1;_5#L3\@1@1b5[0Ka?6\:H+U.;b51Q24.L=Za^7U=5NVP^
6)T;XQM^OYUZE)CcX4O0VcFU[^?g]&c[7ZSDdJ\[NUSbG3#.H3KZ6NF3N[9+<H7F
9.Mc,8e1>D4.\V5HHIHc[G+RHd<eg&E,bdS4,3DgH=gA;B;aI2,OTU1A@D^UR3@G
Sb-#G87MIY5fI@@WT0@0-E-M.->>^UBU8G+Lbf_RR\F)AUR00^Y,645K@/=YT?3M
7?]L1/=WOW=]PAK8Nb>c?8^&-PYbFD/QVb0?:A.->1U01F]K:d2HgMTB.)(&IG_+
0Vc1b68)159Q#])IE6\6(ac<]&)MG^T4AQ#e#H(59,U:WB;@ab2cP3?RdcS>RC,b
)WRc>&W7;[XJ7(^SOR9GZ\=-2]9E?7,.(8ZC1FZM5RM2W5eZ4^W^6K[39POYR/KX
R5S?ZHf#PE.E;K_O:<W8>4:^_WXa?1X&,/R?aEFF0[gO;.dDD47WGFf[6#A[GF.2
+_/ZH\[KM(e\\,BacS4>05#_ZT[]3OAF2#E0_-K@KDHfZW,6-W34J@V,-J=f&2N[
63B5f4DbJ&O\1JVJ=VPQK(#&51=8g3B_4?DTN;7T(//dU\,5cH1]2&[EX]M(VI<U
41DcS<YOLS\f.&_&_Bf4M98?BVDGKAf]b(?L#Z7=Sbg;IQBQ8>ZNP>Rc8X3c3V0+
]X;.@f>EI^QJ_gG^:=aFdAZE-,J@ecZ+R[-=#TZ3Kf+9=JRZ0T81bQQagIX_-C_d
d?:ZZ6&:S9.<]f\.c]<ED5^+<@MdI-#^H6HUBEA?TCag#PW[aD;b1@HHSf0FTWK]
&97@FX=A\_#7&T/d0SJb>Z>?_d#?L&#2=@#76UA68?Gag7,FM29?.LCE[FB&O1-X
F_Bd;61,eH:.cgbTS(\7OARg=fZ49=N)-/7adZ[c_X\ZA;gQT/IUD:\W&f/J[?@A
eRQ-0g5^(&2?JW.=F:gALJ5^_aFTDSSJPd0a4I.FeS+N<3,eQ1O&g4LGBP90;@&G
;E/ML4+6B\SUJKfgR2FU<T4c(,:/X<4eNN\@(Y=_#S4#(A,(>B^T[9.UeV<,a(,6
b3e\2_M^E]Nc^MK[_7\Ab6E03Q@\FYd),c5#^L^2DX@e7cJ27FP-aVM,1(bT+.2D
I<9LS5g0_I#fE;:#E6YP-B1NZJe[N>.cOMPHfbK>Gb>;O^.YfJ=9_1Z_N0IeQSV]
/8+5.]UggKB[.L9481ZWA;e[&+<KKK0EW_ge#7XJKDW7-8VM;V-4cI&a,O.?YGbb
FKCDE]N.dF5HW\)OOBF3#SB+ALCV\3-afVfABER7_JV:G].9^<0MG1-/U,UQL=P@
#6YNbROZ#S,Ad,\8=-1P#<1B.I5eb]+)GBG@ZFdG[NSA250fBe51EJ=8LfO;J06V
d=9G@KDMVL=C;:L)>:^-,eAZV;g?A2(VbXA?I?4gbecUCI9EB)C:6T?DE/1]cMUO
48+AS8(Y0UXLQaCJ+fQ_X\C)I0Lg2\HMQ4#[NdaU]7@c5AGY81/S4-9MH?QXR1D=
.6^<JDH3C0:D-E?DJ>:G^55ZCRB_EK^TU=L4,X;T-)0.\TR/8A3K1c_+g-H.N0U8
9R8R:IB1IU0+RdU&Oef44H8;eGR]e.)QL),;(&Q>dN2Z.X_Fd#=N>UH,;KX1QBaV
A+SE?^GJ@^HK^OR;JXZH;ee,0SG^LANE6F8g&XS4W,^R[;2JaXa/H(L\7Q=fbOJ.
V8NZ()Pf\=PgV,IN@7NFTHJ44L0JZ5AGUd6BBe)VPc]]XE+H/Y]129-X3>BM2B(.
Y(XS<Q6-8ScOO-.?6V,X:QMCZ^\M:10&<((>34:d=EB,1LW\=90SBYJa3+aX_b,_
O=U;>XUQ88P66.]HGNF))Mb-O#?DgBO=Z@H;K89P5,5C.dg4bLf,]1R7XQ.gI)/<
Q,P[-529?W^8+@cQ\[SIR,d:@:WJ@<(YV9&,PD>NDS3CIe7R\S@\@UX/JC\]X;L=
+SXAYAbI-ZMVTV,S72KB7.[K:U<Md&Ud&A;M&+9\G5;a@[c2WYX->B[PdGg8<L<K
^3#,Q:4K45JGU>SCJc?T.:)6D@5?HL4Q1fQWZQDa^@8J5DBRSA+F+B@M[eATbT>N
JN9^;T^bZ(IO=?7NB&-D=6MU<KZ?/S>UYGH.94>#c-K2:,b=(OPEQNR_)#YP2?Z)
TKFT<R0&381&=)#eQ+_abJ<8aU=dCBSP]-)0#L_d867@#UD;0fSOg^V(X,E8?(d:
9]M6TO(OGdE>#RPHLQ#)/a5_]W&5)8=A=+0A5F8(>BJH:SR-S]2G_JH:Tf@\>c98
48V)R-8RDD8,fVV:+_(JI]+SVDJ8,8c3,bV81gA,QRa<VJOO4>P9#9Q.H<0g#aO+
1D^X+.W:?C/VVBX?,7-cD3[R]=OXP_:BWQY69[<LFVE:?@#-b6H9)2OI#:CV)<O4
_&#?a<3PgeVQEZI/8U;CP&]M,1PaQ_[/Z-=L8GH,LT\/:>.gS=5NEf]d>=]D=^]<
=3WUW>B92TW:11X:5WJE;LN.\>5>)Z:HS37;WOJb<NZSUb_Jc<MBX&J]eLH8\UcD
2La(+d_OSLB\M&]Fa<R/I,4;;OA<_NYFZ^M5J]8KWXZYdDV]__/@)Xc@cLQ8626N
N/^C=U3AZaO2)1AH;Lb3d4+-+P@4P=#]I?QQIRe3dWaFW?I99\cfV#/U-[fDXIP_
1KC[?Z@b#)S1V?1JKJYG:U;-OC[cH_M.K+P?>I3ZXE\;d8WO@JX^8+)U]?@#K]H7
\TS\_>Y-R6K1<=Yb0G.d+)/R#O:)YQJc1\bBG1KV>>4W8(N#J)E<<EK?A;+4Rg^N
@^]aC0QURI\(-W/J_7F2TM\89cXTA;(+]1&WJ+-QS=B9X<PH.=IEY[(9F?=4?X8W
?2P=R5bS8^aJ\1ccEQcUX4?(<,&WG]DR+N5X0A+U2KZCA9\Ba/WE>g@DaXX^@+^[
f?9QYL?LfTdL5aO6[N\M#>AND].=@;b4^&<N)_VGTK:9VB=TRUBHP@MD+/_Cb.)Y
]_A,(EQ<b_&QIT19d0XD@@RT3WU4DCQ)L/@[<(?HXFS/?Nb;Q[&GUC_gGfHK1d^:
MXV;458\b,df1-_BbTU3WUa+=EWe2W33FIP((ZNGO4FTU3eN9>65_P9eHYL1YE+F
Q4+8-4795/+K=W/7]3PFC1V6)R=@[L_Q_g)Bd^Q6G2B#=a-e\R?6;)(UV4J\:)<4
VU1<?+M//5#3>]I9HBGS9LYaOW5\C,F=362#;)&]#-0-I)_#JB.GN]FJF-\[ffX)
PGc]b5@M8g(TFRP;7I?846^9)IM@,+L1Z0.KRA]21(9eYPK-;>Z)M@<=@-\@Ta&L
-c^]5Q?M9f7<5aOF;>CRFNH(JBPI[cSc1=<1\_M41O49)=<PYJ8P\ZVL3PReGN?6
0.0N3\<S4C[2EgM]?>]AcfUESO@Ge)MV_dc^/TI3>_aL+NP-C&LOC?,)B;B#8,L8
O;VRA(D5,5Q?V\PKY#>d6CGL(Oe4EJX)(b?-DB:+2\C(gCaU)T9a&@R>EIW+XD=T
UXX2]=cE]XORX8I5DPZSbF5#>G_L;gS(E^a&9>c5N#g)_&9+8LZ(W<&Uf,2/@F^8
^;R\DVJBD:Z9e,2c3e/UKJPbYc\^.a5dWOH)DP]VN=+[4XJe8eNZVG+I5DL)A=-)
J]EJ/>(aZ,EI\Pa>^J:bMZ68eYJ.c+(S].HP3DVQ;1W#c30OB,c,>U^[5FEC99d\
;]<M1=X.23WJ8S0/Tf</D93Q;Z^?O_-:6#(NGL#\>2)/H[e.<LJDJ0a,G<NW88>:
QK\g3K60a8RJ96M:&#E#+J(CO,<bDI-[f/RE?SAM0WKN<ggdIR7)(CaHDE]fV;bg
BDOPWJFK057>);#MQ+9HF)Y,J6,FYW/0\,;4W:?c08MHb\_)3Pa>I]G&7:+H0JR]
>YX>0E6-EPK;8M^4c15T-QUY<A:V?6R7#cF\R&/5Ic<]ENbHaK-S2@^4bBJ&>dGM
)-9-5M_5C&ffR+dC+S;^bgZ:3\HTNOE0#dI0H8F@+:0\efSEI#KU_ReBdQR]EATT
TJDP,OZWM2cfHSK1EB@=WKA?W0O.ZE4EV[DTWY<VV/67f\.^^_K20K]&KGM:==7(
3P8<,RdSTJC,_KWT4\H8J69=C\c;7#P))?;3b.O.P:;XJO)S3M(^?5bbY9-\Ya<A
Z2,gL]E@;/SR+W1,KO\+I0??\8(3@])LLSX1]M_JI>Y&+9A7>.TM7eD1LDK9]6MY
dFe<2UD\LKW=W[U@:+.f9X:d=/^M7F>&Ugf/+96NHb&OV.AG_VW.\#-G30;@PZ0H
.UZg-gB@b\9L.#37IC/F)46J[_AN\G1VX=W=/b?\<VR0UT<O?5QCYL)&:VZF&@4L
:B@-.ANFG>8S7N9AT]J.86ZMND&,0^/Q33S=;UaEK;?e>P1FbS5^>#5LQCcW-PbR
[AH;d6:K&,_G,8IYMV(SVZ?X)KZ@6C;ZaG=&OcE+[(I<gJK7QDGXO,9caD2(e.7&
<J1>H,f?;H5Md=aP_BaK>LH]-^)R.5;.Lg_)S7?@S@LIM59L-LA#F]P))<gOVX-a
Z5cBA<?U+eT:F;4d3GBU^XL<gSdB-Jb.:#b[[6>#_XX=A[<C2-QGSW^J(M#J6-3J
PW:,7GV4TA-RK^?ZN[2I+;=C6LBfUV13N(>L?E,10\<OVNI(P^g2/1T8V9@@TU9Y
cS#1D)K]S[Z(aT.#PAL(=\Hd/O1W5,TSVf[BGf2K1,4+e<N-Tdd@7f>DI#]fI&EV
X6a-Eb937c,CUSE?K6J(21,<K-D659b6XX^RMXH.;2J#]>^_,9]Ob5)E-)0B[bb,
:MBEVg6BL&29:bIE3)W=Ma+##\/2=HR&:DDR=H\EEE&X&X.b?K,e(RC_-9&S8;4M
GG(<N22/O/a,M1CXVY-#GO\R#8(H[MgIW\T7X1EW\Fa=;cQQU38g(DC\fI.A]QAe
S(TbQ5cg6H;>aGQCg_f?_)8S>\bDfXKRQCG#TDQZ/A67(dSUT/0\E9&ZA,[a&&cK
26)d1,@<R-b+NT71T&bf?:A1^Jd.XB5D2X<^Fb<PcG3U3J7X/Y8K[&ec3Tc>5Q:<
,&7.KL9=/LcUR(L3>;dXT55c\>2^.5:&;0feRGGO-fJ5AY_7+8#&GIGH8,[TIMPf
[Y_,,,7B4e.WIJg#6Y&H&2[E(AC=^Uf9;M58@a-KQ#;4cBBg)HL.Z>d<;QS2(.H.
;#]gMASZ2b^\+fKcf6Y;_(:)XU6&39=ecOX&&&8+8MSQccF7c?H3EQI7E]HZ-(:c
5NM4M@OL=D8eMC_],@f:DA:7-GBX4gg^P#dH0Q]FNQfM3(956b>JI;IfM6(7BJ#a
3)9CVI@dY\&g=MI;AbCJ7T1.eBgA)#K?<LH#2;aY0FY>b[9cZILY</+PN\V&[g8H
T]>O.?5Qg8&(W;&c81JQH^D0b,g9\&UF+N;VHE/USOf@1M@3d18E\;ZDYEC6-3dZ
WBR8deVI-BVI;45YB<Y;L#cSKKYK/_f-a?=_SHbS-IeQfI:HPL;>YfGR,SJ?K1D&
+M4&SgLMZ>\8S-J]1-W\G(1=7K\@^QRUa3O0E4OX3FZD4aIc,AC;e<^87f?dU;ZA
S3eY=?RgZ]S_A.JYdP^NO@9ZcDXRP544FSfWK8aOGf4gK@(?YFW2gd>bbLL[+XQc
;fa4<G^K[>-e5T&;>R#VC-X?=Xe]fA3PgLH<GH\SR]C?8SSLZDM;Z?#ZF_#R<WP3
QW@YU>#>dAd5/\Q/XO#5M.aT\Acd6O?@7G2^SPNOfA5?:\]7Tf[Q=4W()5Cb(447
0LI4&0,4#FZQDSC,A[Ca?9a-/1TPQ:R]@6<M7SMHJ=:X11f>=df?eOW8LOP=6c1<
BVH+Q?QE=HPE.c17BW1;=F#KF/Z9A533AFPXOV.PU.\FDCC0G0K]XI?T@-LMB3GX
(ceY8/b4<^U#HKQfb;aH0M7)+FT__,c?BaB#RILIH]^-5e@c_UL&[?Y#WK5Ff@]B
VQ/:eG)O;TE,<dK1R@L7-_L4J+;J,DAD;V;_2Z((DUT_9FJLa1c@Z8[#c;L#<GE;
\[1gX^ZG0cU]F3J:QVB38ZM5-H._UO?I9]KD.CRRe7<_I;V+IG_]QEDT_BF>fM09
^@8Ce[;>(RZ?G.F^4+#&J:#P1Zd+@YMH5@]F;d_]OM5c/Cg7]>(#4\N8_T#VEgR2
[PUEZZ1gN1T_HSd8GPMZ?[gU^d8e,)5YLA@7aJB/]Y[BSE46D.,BaAJ//\,[QK#^
a:8/@D]#S9;@;H1J4#d;?HN2D0@YD[]@RcdA/<A17J=::dNEQHG80O)fQ:F#PD6d
Y6#K:X#R&AeLW,:1,7Jd&79]&@1#HUI?.#7aZeGP6Y5YCUBTKS;5a7H<,V1NFJP:
U=@-dH=fF1V?OSHH18@d]<3EMgP#=:MH[,9/>[fd@_7=A9_>/KWdK2&F7>6WAc@\
?>;?eP06).3XM5<D]TSbG5Yg-:#OUWN#QP?f+9,DTb5(ZQ]<cB;:7cJEE^aeCW12
f5O>JFN;L4[9U/8-g&=Z75+d3.24J6_d+OEf5g>Ug8Y=Y=D^^7#C\<-[M5U8+e#1
63VD_E)SM[B[5M723)]1D]7B8eM8IBI=Ga>WM15_/;T6dX,AK?U#bWYQc_B+@\V+
QKFBeU38gG?a@#XWXNdaNde\gM>:/a<)^P)5I#T:^H,,_S^;M?A9V)ab9S[RTFeY
dK?#]VG04FOE(dRTJ]LIM[TVQWR,GOHK/J]C0aAWbRL.BDZK14Xd8]8eI>+N4?5(
L+=]_QfRCC6,AHe8HD5VW-SZFd^3QZ>9B\TAU5DE]P()LL;&5/(cTc4HS-fB:CSD
\#[):.XIX<a=,/OK[EQF53#NeZe6P433^^V^:SF(,^aHQ]P:4eE&[=(Y.2Y9^3?5
.cY)CN9Y7SLM3EAHXd@\5GC)L^.XGC^fK:^_\FIFSR^<<=[S,W1ZQU3Q;LBY7Pc2
.\(2f],f8e<PA+0c;J5gBN5aN#Z\]fQQURY@BROU8AeDQ5@/ZA8W:PH+=BG;4Le9
13>XUeb1G?2a+PfP+B>-/?QGKd/D=/H#Cg.+KHeHH#XU#/>bS[gEX[ZFd#6\0//A
V9-@-_dcP+ABG\T+=CVOKe0g@HP[,>&8IH3,.A;,-6T&LgOcb##J)T#^3?U<eO?T
_7Q1IODfSL2R^b56/Bc_da:CJ]23YG;ee#-c)57gGGf#LGX:I[Z1?VQ614_6CMM]
=Kd=?gOR5QX<KRZSAS.:F5J2,18=MDDL-fN+U09IL:\bg)9e#J9&KJBMIF;C<3=B
W142\&@(-gXA^FF[daW7Be.fg)ZdbMf[^/7]XLQ.UEOJ@93RXM#94=D8=>BW7B>(
g.P1L1c=)7bF@WM5d?/\TR;>YOR&D7Z@1C,&b+4c1O#[^4\P6D5F>+=8.CBL,@=T
0UUeHM+9d38-BaP#9S=CCg/MHbB4HH;Z@](L?MYaV4(T+Q]\):d1<HK[ZJ+X\_aZ
QfUL)(\)D4:DMcRMK[FZ:15cPc3aCW1&>G4(Z3+8?ZNA&dR\]cJVFdK2;2SQSL?A
AIfKESg-[<TPa>^3bT2^/<f\UBO7P\PSUF\K-F1L2QQg7=]6SN>[STOf+I\EQ&gQ
K3QG2X4F:POW6M.\dVP1,392S<KN,V:fLA3\>5eSO8Z9U;&2#.ZH?3O2R:,fV)P/
#0GO:VED;ODGHIRO#(2)&Q3b-QJ\)Kac;)Jb1+/^S#A\8IbFZ;1<3<(dJT&U?_\a
0C^?GKO4F:G=E4Q[F^Nd5BD9e13F\ZegQ7?\Zd5d2TI&;;,ZaPQ@>C-5B1562Z\T
^[9fCT9>_YZ10HEE.gd]:^aZ@E<,RJAZ>Y/VZJ@CD]+ZEX(g+aG.G1.\_e+aFE3X
S_AEb@/dCA;^/AUKM\#V0T8C7d1C7ZKWM4-JV=.66\b0[B>Ce=&4+:cNU\+VE79_
>7MUSK8PKa4;-AZ:.CFeA?fF9+0F^2CY.\7OYIUX\Z,53>QY2M)W5^2\152OP;,B
)<T2PbL&NCdXS9#:_c6)0W[8Pg[U^0(-=-X+K+H3[[6\GPdU-/b1Q];b.SM.J]Z\
K#2ISO(;PF-,+3JA51EK1ERI/WNTa6[S5MTQfUOB/@#Z9XW_eHXEITG(()(4LWcS
\.X0B#0V60dgJ-Le4:<ZPHCD7..I-0TEF/ZGN5Xb4.LVcWV2<e70)(WbQSE-([,O
HB#S6;9_9f_C+I+H:Z8f1RCP5bS5d.O227#@=Y-KBNOE#38W0?F@A?JB)e5PP3@0
W[=EBNPfR1eRVW0#)V_H.M;&#OB5#>a\U9R9S.B,4H2dN<3+Z5;ge1JfN;ZY18F1
fKWF7b\)e3ZgUV1PU\YLf[BV],fKf6cc6;R3Re)\[HcW)dMLJ)6,GL)MWO-TJV^c
fWW+FZ:fJ19(Q0:g_dU^#f2\]/CLa6X7AB#N]Ge=g#_6C.1047)6g?_Tb<gY/D;3
HS\Td2V(ZEY=2-9X=?24SLZ9PJ)8-BAT?ENUQNROB9R6P31I@gPK^B]b32.8ODCQ
bIX_)g<N+43g:,cA4XG:T,TFPY)J\T5B0P-I3c_gG=7.:^&75JEY+f#^65@B@cF&
bK6\^YK(C(5CL@QBI1H(NMWI=M+=WNIA8bX]-aZ-LIWU[CH]2^7&J?G:61\PHH;9
&d7e.I/G-3VJf7O@:?8/Uf@5;8&VQ]&(GgL]I7WJDQK;f&=\K@P>=?T[:<:BDAY)
:F1NBb?-&d6UZ>\Nb9P@L@Z&[#I/b/Q\K,0UO<.2K)RI>>[:XEd2B^=9fSe#6feE
)+>[Z)11X\W0JUH-?KIFEI<?PVb_]g#BbG_GLBJ(2]PSEaW5Z&R]2?QH9;Ac2(1P
/9\9aa#Y#5WUKNAK<,3^/ZT:+\4=&ZbR@2<F_ce>>QVLN4=7->=(I>Y1F6;^TR&@
E;3T/(85=GEMaRcF54I?[/WH#P:Z78D#a:.Tf3:c2VZP/d):L#C[JWO99<(bC>0O
JF]P+:(>CGC1CC#W:>;MZ-S9\R/X?J>J3JcXBUO&TO),2=E[g@]H4.ODAK5;^:ZS
8f3a\KSC]DJ>1XedY_XZC5&:7b^-gH[YJL-7ef=5,de)OWY47MbC<(]KMP06.eE+
7K+>OKR#X(RJ8G-3,-cRK,9dI<[;cFEb@Y1BbUHR<1>b0TNHQWKHg]^&R_+:<N8A
3NAS\N8N(<PRWD_-?\e/>CeYI]DGQT+\B&01&ab&[&T4#T+1NDJPMS#LR38/8OGd
C765ER=)^9LRPY][<EcTCOC(e47FF#/(4bB,:]]P#@A<bX4OEFcJHKcV(7_4E:H3
^O0GSgVgR)@>:2c?3&5N/&<F7E+B+3?^@-U;4R8WOS&dA7#V311+O?IK^3.D<7S_
]8QUF,+8PIS;]&63W,a73APO0e1@ET)&JF)J0YfY>GH9HbBIZ:D]^2:=GJbJ86T8
2B03C[6[K0Tc1-_9P?0J:@Q\2:acf3gP8NGgT28Z,TK+5QN#(&QR=WMS,1XB9D3V
84a11GCe_BGdZ_0WdSQ)g]T;8:^2S1SO+0Ac>MBZS\@A@[K/ffO4[CQ[SKZJ&QB]
8D.,15;0RI&IL?b;.J0O5F^:@:?#bHP]H>V<];SOG\:EN/(8&)[UaEJd/V8X1P&#
^67?\D(3Mf&5#,/54dLS[8)4f28df4gH[J0?WA36;4107G\KL[W\M8b1VNP1Z>S0
1YM4>DJf0MK9aE#7FSAf:<I;-EXG(S0f)G<BbeIVZ#\Ccb_\UV:L2X;ZG(dPO(c,
+,5]AP<[@RF<>[MPA(F\ce)9.+3+[<P-LU>Y<9KBGH_+QfFRF.WfVVGJe^-HJ&U(
eS@S_CDCB[DUT)\]6IHQg-X-7LbA9#[2=PeDQ(3Aa66Q[5ES5+.E:b.TCQ=@YcTL
;KEH?+L8HC@[B=ORR&PB\4fa9#d[@D#CD5ggUa09+-[\cLd(9<V/&\:]U3^b<WaJ
_B<[?>ZfDL.>D^eA:TZ1E-?6H)f]0LNJ22[D9K\<)?E/be4\/)VaINe5]\E3S]-]
MV[1H^V\,MPR\UQGZH\cf>X/&+dIe;0PGLFTI:NOd;@gD00.HVbETMNYg#Qd]CDD
569f<RAa1BD=8\N8H>8:ec\-5aWL4/E8)YZ4#aNE,bI1dYGSVX10NQ?OM)7P++&P
[)ggXg^-N.1e_KMZJ/gV#DKgPF1D_E9[IO^6^eE/R64g]:T=gQ3.PR-5J,V7<Z+6
:B@E36R9CIJ1gZ?J=KA&Qd1DDEK4KULALg>eQccSY:@3IO/2aSTP^#S)gXW]_K#S
.<=6+b?f6:(dAOMG5?UK-HDYN[/Bd>dKVLY=-0U\gfM&DRI_a-f8[/c6+OYV2.6S
[:2(Nd,BgAXT30]=(+?XPf,e&S),JF]-7^:JT[O/S/0bF&,b[SU8K45O6\P.17;)
[]>TN<.UNTHgOa_,0c5<#[A?e3C&a4\HI+MI_.gCf]FUJ-:JI163CFOSc2HWQWWN
3WaTK[^/@AgN6dL+8;5Jg_6Q3-3-fOZ:2@O6Y_I28XDd;V0^#W+U)K4LA4e_\U?R
([6GE,3B>^DU;cGXJ6\A4^/<>d;Y\\0UP&3:9DPSCV=7G0-U1&CcO,?X\<]dPVe@
.>ZXAcT[Gb=;BYS-E8^Ob4>DD(Cd<,<..QbD@Ra;1<Y=<XIBZQNL&DOF.U&/D/XF
@?;\F)OY_WZ8&(XQR0B-MLWJF]VH7W:aIKHVY&E=?M]f^Oc_g_<O2Z-T3d<<L_U3
=(bJZQNY;<1Df>8,89(Z_=2gIE+cAAXF6)BbVK[E-b^2UZKd:77;KBDEN2IM\S/@
O]4LCX8>_/S8,BHN9;fE65O^?2>:+T3_W7\f#IC<MWU.<(7D,gU+0N(]/H870>&N
U36@C?IG..CY())\=5fQS(3_-<EAT,2E:NZ?GIbRR75H6WbPOIXFXOQY,P-ea@.;
&<QXPA(E.?c_R.gX1X1)+&QM4\KKDITCQ[1cZa;1?&4(bBO_?L?4[CK,NXB/Cc)d
N,gZ,1WM/;dLTcbAH4X(<S/_]Je7HDDDD]LV8?LYC>JC&S:PeL_5,WM:?deH)5Ab
X7P>dV)@Sc6WZ/:&@]d?S2=eE)HD6GN;@^F0^@OgCD,6L0R-N^a2fPSb#J?/L-J6
51UdY?=E<gWK6__J]JCP&eZR.GR1:gAXZW]T\.4cS;\)IfLQQa4:GN8U7OHeVNY7
bKb+4MbUOQ\H<&c6=]4YTI9LHC=K3A@.\/7,f/IM35PBM\Mg]F,#>@C.;/H5-CNH
RQRPDa(8(adTbS\J-A_Ca4=HE,KZ1.TBc(#:8SF21WCgc&9.dSQVK?63e:)eP;YG
<63a#eC<Q=G(:RT\37,5_aZ\QT[:L<?NeMP)&^#KY><g,EgGASD<1b_58NU,@V+>
?^]P#]W]H@6BWCGUU6=SI:bC0D.S9eXU]T43eR_^+fN]5+a+dP_\D5B]?E9:#cW>
3eMDFFIc>IOM:,Q^faMO/HRVH)>.9Tg99L.M?Od<\7-,XCaa7KEA^.dJ,g(T-),&
dF=S&Y_;NdZ#S[W,]dc\A>[V:V??H9[BTJ>49KbXSZM#RDc3-[UPM3SgcC@AO=BI
gF77,FE(#2;KS<7ML&/1AG120]^cd9A#cQ=F0/bXLUcW-QJ&IQ@YP]a(fFCH1Z:f
[7/Y+b.d;)5I-QT^00NZ3S:LT+JfG(J:>gAME1^/d#-8cTM_,JECK0)-UC.<TZN,
)[D8/VS=<d1Yg11JV^8V]/Aa#L3RD;S\g;Q3[/(D3:K\1aGX1#<BT/2M&3@Z0V:E
b&GS/H5D_K<54VW5U\KJ)D(#D/dN\eS70f)II^QM9=(,KgdMD1^HVY;\)\;_U?If
8^LMgb:3MCH@1:Nf,)UWRNZAK^&YA>d?\IaafJ<?<.L^&U+O?<XSK]SaIEBZNWR[
YTK+H(1ND,//S[[W-4]PGE&d2KTB2J<I1,140K)G[bcJDebH-[T0f(9.9G(.6&ZL
D?M71UFA<:<XQM1W.E3@]V3S1AKSJbK9aX??>S(f,-gCO#9@P>]@P:_gRJL^PW+/
eBZ2OH2XAMRFd^HeU_Fa3QP3fdL=bU0AYRF8gFJ>CL;Og.B:d)_2WG_BgMf1&b&&
AYQ#Z7YF:KI[^-NP6,8XK?@/.A5Y?R+d[IHgZEd-4(?UTgEYKL7I:-=He:+3-U8C
5W8,AX<MF,N]T\H\7>1.L^PP?OY5a._4D/eJe3]TZWH2:(9\+6>:IY-05_ZS;K:]
]M]XX-?(FKZJ_W:5T01SZ)@AIBWO3Y7(5&O;?NQC=<R5F]TG>Q4JbE;4XaSW-_L4
\E?[VSBDFCO+I5/9FR6QNNZ-82=gJVeFE_#97+^2YYC[g1+O<PI6c(0,LVJ,+?/8
9NQNWL.R>AHHdQAHBdH>/Q@S7dFT0MZK[.\Q/84COXS9DTTU-K^3.7B.JF\_9ZGU
\Ka=f&D]gcB-BYF,0a9[d2MN.[>KN9JAJER>-.8][D\+(e@B:#P-e39PL=Q04cc0
CdPE-Q^5g1E^C8FO+&QLB3>#\FOZ;Xf99ac#6)T=;&X0.e;5gH99?B1<-FXQ^(DU
F>#JW)eQJNWMNe3^2=W=#I:AM91B9C3Vd138fE/Hf+S3-Q/F#_C#;DB(<C7>2DD1
PQOXH]ACO;5f?WN\SHZQ?)FZ/cA:0?8Ia/]WS#_67D0KA5>6RUD9=L-@\AK24R_6
@M>216[]_&[KRfe.M34T60VZ)dWRcONTI+Z)[4EeEQHTL6OSP)-<4,C3665#HUQS
(HHe+I+MKc9g;SV][KbQH>5d?e2LF^8\=^JP;WT3>40)&8f0aa9,-ZZ@CF:Z2E:U
3#Kb9(J^bUN=BGGAVa&XX\]g?O4Ic0<>)\R\Nc__b30a_^/,]?_NN:3O059B,<ac
-fW/6WNfI:e&XbAVJZ_M_ebYaF+6]0X>@I1YNQPE8&.PGI5:7&^;K)68(X>9H6GW
R_Ye=BXH(?D=&cF]<^CFA?eJ<Z@)2(9WbXE(,aIORDaMV.W1\46H<FQW:/AQ8_R0
W(TX8\bF<9MIY9T:P&<W3]d]?Je\R]aH55<@LEaB9+@_LONQL9C-JRH.11FRQ:LH
-J\N,+ZY45KIcRI[<51\6+XZ2/].L79a<0,AbBOJR#YE74\^96B8c5fJI0<+2Kc@
-0\3YQEd9.NXB8;OEL6B2^6H)0d50QX8;Z5b:C#6GI;eOILA2DQTHX>IO@O+57d8
GAaL2RWBQ:2/?V9BI93SE)?TNE(_Q;#&&(+_YC2LQdP#^EW1DJe1/:HaV\-XZAcC
&I;c27E-41@cV1UO>64_;,KF.e05K0cAb6?4-9g3N^T0R1B2DUa:@9d[-V1P\604
#>a3VT7V<N+[bfa:aF6T\75#MXa=4+P/(fSD-8OW>5,>F[M;R8+dGO;JXGf/T#VK
O]Q0=PX;VJVXe4e&FI;P75[]#&Q:,Ec9g=Q]]#KC]-^KLfEcd@D\1U7H]#gHGJ>b
^Q^FDORXH4.KUR0(^ZO<PQ&-X+)P9.C6P4ON#5F.XK,N;@?b1\,+5YcQ3S7J?K<4
._11QC6#[1f@?EF,AF::46Q_2?6Ab.<I;36@<3TOZ),7O4T:54CTR2<#-+DMf4=Y
HQ-d5NJU.Cg?;d?\Ae]1+8,=D;169?:9DH-.\@&.9[#IS]\[(I4)GTO59Y2?KU0d
W/PeH-e@GEHJ->[HP;FTB^_\aMb;IRH:OBP6\Vaa)MdUWd_IbYSSM26e3[c)6,8)
Y>0AT>7OPTG:O>ZUegZd@_8UAL[\,S,@:Ie,ZH@@=N1O+7TR,:g0NE?,ZAeeY1_/
eb94QReP)S/:>PN;W^+JF\[&bJ.;cT7S/3+Z18WgXa61]?:LIScB5,#LB]b[BXFH
\4B^1:f\#GY)+9AT9(UIE_SM@C]e_.7HU+6M(?N>H0G?cd@c6XE84#ZP4B//8IHF
e<e5XbOg).@1gB]<K==YbQS1eOf_MLAR\fH#UBWB91XG<K\?.P;aZ\=GdVWL;SR:
.LP5aYD9^fH=dPMa2^5I?<>S21#RVUfd8dgc1YFM-g>6.,BUNV<;/Z#FJ3gXCeD_
#cg42Q(:8O]L9=d30f5T,2PDeeN5Q0fA=AMC\>C8R=6W&97N5U>@IDM29)3YD(F@
c[\;8/U=(;4,&I9L;N;Kd7JKFb.HI:G\b&F,PFcW,-2AR>8:[bgd7DD594K,6C@a
+3DYV,YcNUe@P0,<]>TVDb-[g_([YL^dV2V^OJ<V:X.=I-FP.T,fT3K6,58O?QJY
.Y.PeBccO\,e,#=0+OO:(?BfW#6GGDL,:<?]X(GfH#-4Sa[>dB=;FfeebfeXa].=
+F04e<;\-5IT^+1MU[<[.?W8_eY36F/7W<TCI4NfE]#dMR6[G2,#^I8M.W,.NcaN
\P]G,gU0TQ#IM5C=6;4GM#[T]YKO/d7_,Q@Gfc=\cRF,333f39)JMJBNT/OJa8<d
L]@9VQAJB&_O5O6cD5[=DNXI@A/(Rg=fIQ\g)[Z;ge2NDZU,_B?AMC9MfSEaN[;>
6KVKOD1^&/8>_,O3;<9J]8G6Cb]B>^bI5?P4;]TcDA0MWHRM__<2?0Y<U_De&,\J
Dd+J@,VGJ&DNbV=C1gIN+T)(;:8+E+)bAZ/1:?0:3OZceH,UM0-1+H71C<.;&YM^
:Fg(\G=2Z@e^#PP?VFbR@2#c+_W<fQO<CZ&W1;RdL;@59KId4f+U]VS(c+\=U9MQ
\A<BH);E,cI)B8[:Q_B=_8W.VbcX:8I;;[3g0FA0_/8a2a^\+1AL/g6YTaf]d9K3
TKD_83-\cRM6VLY0K[/eU]]E-?HR_@N>#=X4G:@-)O.MRTMfKEX,[Ca);Fgb)fG3
RfT[(e<XcgBDD.5(I(>::.ICT:BCKH1D8g^N9ORd_dceIc8d;]5+P1?f3Q@AP,QN
Z,-^OZ0)NOQP;?^eFc@OC_](0/S/e&0Ha<SPCa4IPFD]@28VfGRD-XfbQZIMO#-K
FdB6ef:g,e=N8K-KbWK@2]V^.6I;PBL1P[2],^T4=A/EU?VURX(@.9G=-(Z)T\f;
:CI6#M>5N5N_X2+M8+OfI<]W>b^=\[6;a#0<c2Z1RMFCI\bF)M7?\8DDNATZ\Q+1
0_b/F\HPg^<AY@/F0V>a:U,[4Z7:&:3W?WOTV/FS<7d#2&HXI_.+IR/6J9eOLeUf
@2OV78P+@3H1^;7NF/SBW:C,7T@OWMY.7,d]])NJE41aSN\WWS_.0e.\H?CNaE#[
R/9?MD<?.3eO27e?+&-5^5Ve&BY+WT]C65,U_L@L;;,f0VP9=MQE9VaN>[]K1;).
F2UO\([<XLA5Oa0MOBA@0R1,(FTRZ(dPf3b,c<cN\GTfcSXIY?R[SdM6D27KZIEA
FeO,=KCONS-S47X0[98,2GY:+AFe5]-)])?/YTcJLF8MOg1)F4E/5#CB9XU+/5[G
Nb7<U2XJ6+KZFJQ<N.(aI-&)3(Ne(IEa=J(SU),/@=^@4Eg,GQ7cDcfMP&&+:RNc
Kc7LYd9@LdCKR]B8CA@Be26R--C()/EfCd=@8^6G..:RR:KJCC\:CIa44,,I)dV=
U8/YV:dV:NVBdTY752/CNG@6&d[Q69H6Z1/17S&)3:_2Y]0Pc_fIK^X4Pc&9@0F5
OMabCN6+]6S);fKc38>ZHAN>#Qb^1WeM047I64bH[Z#_NA,[Sg;3U0[B.f\Sd#@,
4:)gNP1CXeQ2f&5#PL5O.W=<6H6.=dKC2N=FMA7-(3c&542_GMRT;^KF#)KTD650
E[5f:W:X.&T2+<(?K3[CH,O5H=I,)I59[/T_cDL]Q@I4g\f1@eL.dAZ)O25-?Ga7
-TJNQB(_M.+;1W:\(#\PK>O>K?KBLUSE4]8:P@E[<S/gL[VO4.H(>57Rf1?D439F
X7dCg&D7dKg>KCd0-IEJ.Aa14GNb3#S<8_2UcNeNOA&>P7M\Z@d834c1e&80=5A=
6=Q#E=YPb\LG-GI.1,]/@bT7b^1S:#6/d#W&[@;#7d95b/S:T<9b69W4b9C<1W,8
MIT5P9KD5I\XYB^3)7UNE_]eA5fGRcDTZ/W8MY?e:2DELc7A:HL22E).Y+L;C=87
ge:7bH9EL;<AgQKK=F92#:aZ3;Y6]+@EU7.ZIMCaDc4#0;UcE;ZTXZ]fJ8U:EB1A
Z[6TMJ<bM/PMN_@147S8P@c-)_Y2@@>bG[;Hd7WQCOIEd+T)M/[\<[gEIBFMI:3:
fL(e#\9XWQUb)S:M.7cJ@>UE/a(_L0CIHVC]P]bTf)/)FTW&G&<(9A\C+[YH9)(<
=?I&VHSW)8>VfT3V^?QgRC]@Ibb??dN2O0eKE5>JJ0E>&V:2NZcaK_gR/0.)^0+Z
PW3ZQ@6<L7A@UF,669K<8T3R#5-FA\F.8])8>(5O;A[bT4S&++&I10_LS_;R2d=J
;a>>@^7;DVGA0f@PJ/@ZACZ_ZT:F_ETOK:QfN/IaM;F:TX8_>g2,/#E+Cg\]-Md_
Df5LgTO7I):B&#6OM&:I1^U.KFddGC4\[WEZIG,EcW#^NK080#D^N=A1GW@)WK0>
PcX,_G+:-a#?,:N[#3HSJIIWg>^K#1ZA;-F_S[:(d:CQ0K44e?(_)V.HK:?9/?F(
;I&2B:g/9#LAY8:#RCX3&\>K.Va)2PPCE5A1P>a[X9f.\ON3;.Eg=bRJdP&TMaM[
fc)^de?SRR[\?e7c]C+=GaaR19b/3^/c>3f:SgD<@>gXgdQJfD+#+(cB]D=(R(4P
2SS0P+8+5MUE@_^K^^\&3[U0>:GB-D0B^K48N0b_DTT.dU:geCCZQ;[dF61TF&?#
@)\Y\8da99;@:1U4Cca3:b-R9238acQ/,DFG6S:R2^M;GVb^:-<HdH\e/d@3(Gdf
XPSC8,HeN+-e1fIDfVW5V44EAZ2W<0H+/<4X-,0fdXUL/-]]RWH53&:?aL-,4R3Y
AB0JTTb]bCb&a32H<B-7RN-9U+b];gG0>eI,C95P17fSE7_4#,aJ/0N&].d[<DV&
NEP-#_.HQGbbc5IB;>+],FIaG5\@b\7:X3/O;D@1.B<<=-RdR[Q=FBHZ<Y71([e#
DI5WcLR5P9C(GH63GV8[fS&T[VbV2ZOX-&e8M=9bd#/Ig/@0/FUgc_\E3.eY61)_
Xe4eF47AMI5T[;_TMgTV77O#)YCKE_U.)?+6SC;#--ZE/UQ;U53BWX=5K5UGN\&P
\^+=Z[)_cD)UT+g]:X_7NP3;P08f)&<E8a.P^g=:HQ[8A.W8TGX:+A+(Mf-?c:NM
29Og,KX=&dC[=;SZ3P_6YggdC,+-0LUP2,1Y23WcVa46_4DV5C/\OUY.;/E8dC20
?4^UV&M74HS>eVgKT1c&@afW=VDL_aWNLC-AY1CSeOcd=E<CZ:Fbfd7bf>WNF#<Z
XT5K?=a^MagI[B(fK9+_UH^@EfgQT)[ZC29;0M+J1FdPX<4T>3T-\BX)&\0H^\0T
a)<ZX&[NR,d?GPWP24(Y_M(=a155d5_SAM2&8UVB[BPT(UOVT&XVdH3ada)>A<<S
L5]cB?GTT[bBF-4,\HHF+N7@Zb&[<@,@Z0?4d461+dbc6&E<JL1G0XFAEUdV.><3
ZKOFeG3,Y_+@RQR?#fU0J5O\3(+9]&L,\b][H&?01KHO:BbP8-NN:]F4@Y,WgUb[
2TT<YH/2>e2=]_A?EVDP,?AA>+_BG[A+62?QWJQAF.gZ60R96BCQF:@e\+>EYQZX
(RE0-;cAIHZ0D(4>5NX+J[55A,;edA6TC)\P.-7KQT3OH3QeX9DPAWPe0^WeZ--R
fKeGC/P^U9@&\DII]LX2#LT.#dA1D@:8c3H^=(>PJH/EaBFRW]-H7FdMg)PDUGCC
ZQG&W(HIBg9f2;LbRQb?RB(PHWf[f\e13.[4JF<=>T2P<+.Z5TbCe+J_W?dL/0#Y
29B.8VBdRKO3^DKEKPCC1;PI/@<62549-G4\SFPZcX1LLg@9.<YQ@]=IL0ad]+=_
1(\YVWU8>Q7d:037P+Wf/G4KVL@JYOTffF_0QZf6=@6(N<G?@2c)WO&ZN44PS;)2
S\]9R46bG8ff\a9cPFV][0OPe0.[[41S.[D<ID0H\O5T4I.=RS_EGX]/]?H8ELXV
MB@OL@_:N-R:S:9fVfa7X2K2=O_KHV7PS#J5NKbK?PA]/bdNHN?g8[RW=(L@YDZa
V^?S7a=bZ@cHeEQ/_/.O\[V.-=I?(:fSM7ALB/U4(CWYT#,_ZX7e.VW^2>ZX[BSb
1c.[MD[5GZZ).20_1=g2KKV7@^Ke..de+V+f-HN<V_G/XDK-a4QVa>C&TNQ3O:FP
b)HD[,:K@_gEg#dRODc]</JH5g.,<0V;e34:[eg=Fg)?DR:g5[=-1-Ec3^6F/b+P
6BcUQ6E:(cD=4.GTGZT=2CU+BVH?O5SL06aI,=e)7dNXGa<M6&Z9<:FCK1bK-DC^
c-(QF@bU2>^+CH2:(0VS3F^)C,AdD3>)eH?7U9=TB\f#dSH]X+K3W,f7TNLD,Gg@
]JKgD8D,49a^B<A]WJUA[a^@fHKHIC?[cL-DJBf6^ggX;_;?#f9E>IHJ,0c?05NY
T9,dD_8,=_b<b25BeA1.HGO7/&P;2;&7:)U?M#M==4ELe79[E;U3Mfb\;4N.^47+
.5_X<Sd<I.(RLY4GTBc@cX\MVeJMI+_gZ.AJ=VJ<I<UBQ7MKTX_C^_/#CX9fI7L&
=b7M[S0H,4AFL;+6W:O[QZXW>IIT\Jf?O:XWG9d)3g5JPW9(\H?5H:G-:ZMU@T57
H,L<Z5J).7W=EMCJR(QSEKaP@DFg?ZSHP8-&?K25GN#cQ2>R=[VWggUZ49:BRf3K
(8(bYb)H8+ED3&U_?9=]7B4AV;T,#:SDI2b?TMXcTF:-5/[F@#P#PI0]HCSB.IB/
2\CO;U)c-2LM(fT,:(UW5VQS2,EF-T<YGWIZ)<Z]0RL5#2+?U?6K89ebO__[1,/c
72+G]9M<CXdXe2S)_#TJ,YBOFGK1a:gebQ>AX+GRS_Ye:c.d6;T7<<O_?ISX\N6#
N\O5@)Hf?X/#=Zb(PHOC4^FI(b+(PTFe+X8EMQ:3:VW(NZBXY,_I.NG^C8<(KVb7
3@8VC/#83aO+cZ3Oe46+H1OYJ^Q39D1cKVX@ZQ>9HNKdRB]]\\(Xa-11ZH5\]+1D
RfJfY2_9X>cB8AdeEe=B9gf;O^#(Z_E6b^Q_&AYSH32BbH^X4+6K.1S2dEI=e^Ud
a[<OfJWP>eUf33Zd^VK(1)C7K^HZT4RZ/G+CNP1NQ&Y])Y[2b24>VSH1g-R(>4?Q
LB9fSIe,AFVOd<1[DGS[U273fDL7I<UJW#0WMQAI[VXXL_cTL@CCPQEN:E)9dO:f
.H;G@MY+UW>FZeRSVRdNVTAO[HLWc#3)<J6f[?YR/9NTf9-?0NSg(+1bGQ2<F54W
A<aWg@\>>6IefbfBH0XCLeEd1.4B:J\)AcKB/b]#\MYBd^:IKGR(GRaP/eVW4^<7
DTS5dTWRW4R+1XSY7[<aBBf>^1;d#+\<O:H.V@]])]G6,]\48g@YZZd>c)?E]XdN
T9P0[WR2F:bQ/?f9M=OV+]I<BA(e<9-/d=W7YV9JLY9a#ULeV56YJ[<@GOX\Re=^
S::DX\G:^=0I,@@fZ:_WgC>EP_[=4KfK39>E?VDL\DYOOBZ.32^D4J9\/MB\GGX:
dZTOfO6@AJ-;ZGGOSbK/#A^^RV)Y.0R;XKA3<_NFD&3?9A(K07^/QLa;-T7Wa5IS
M-B/TB=,:IV8564=J0RR3=<NBRCXc8+0B\&DTFRZ:fFC7ff1bbT0>W,R?HL9XZ4)
OA4eQC8XD^^7..).6D)=LI68HHQcZ5eI4HQb=48H3/.[<Y><AFe2>;S4e1^=NPA1
.e7fcXNCV^&T\0H,Iag;/gD:e\\I.B.gL(U6fP#N>SS#Y)_8M:MKdH_HBMG6_?M:
aZYOP?24OEb58c32U(Q,5#HQMZ7=10_dD,27F]VFC_gYN[<?8B+PFJg0a&(TH]Z)
<K>#7NLK<;eM;UbGbTa2[U3S_:NC#bY;N5./8T1;@0[KC2=-LXc)_52b:AJN5DWd
(<c/(4@6G(M:Xf3BP&>=.WMT4c_SaI[+C52]3LVc:@=R>fTIL3-SGVb]KOa0PZb2
c^10-b3[6TaJ]>LX2>-XdFKL_Ec+NGTTCK@#6_f#@R-5->4FZPH&HI#[-<,]YXMA
\Y_KOX0<M_;L&:f6?G\584T9@=WeJ1XYYWFFc)862D:M-)d#gg8S+O&VR9X=WU)J
+b9JO0gb]=K:3(EKD[2WN8=BC4>aUOBTD/5V.@U9MPf_+:,Y@1IR96_40GQX>Y@/
7NdNP)[HX1X+bX78\Q[WD^TXc8a)a(UDEFOaFMC1U<F^Z4XF5#Tc^94;MbU2T^C-
.CfI3c6gcG>Q4T<H5#U=8?NNINC=,0Saa(=KKBYGJK</E;dX,J0,1bR-\3Z>2F2d
Y]3P^?af.bPCg@Q3EU/_+.gV:9ZJe:Nb=O?<8BK/DL^(#:Z5e9US77bUM9([GDJY
G\&8&4]@Xb\6NEEdW4;&7JQ>g<\YC2A+=H[:APc0LYda;eF_89C2N<;V6WGef#g[
S2/dZ2AUZ-66SeDM>96a9QTDZTKR;f6>=TN86Z(N09RK=@gPWaP[Y@EJ@5[VN1#+
SbTT3GFb]eDQf21fKX^Z:Q?J[/fB8\6ZEHFM?RASK864fdUPb>EMA;/0#D3&9?dP
N+cC,F2MeD9US?NO8Fa=Y;,HJge)LU.)]>U60#9]W29c]ZAA5USO;+gN?[-+#e6K
09aeO2:[R?NOK<U5WeZ(Td7)Dg/(3SFPa>fQ??:\^IVR<H^BV)DP_O9g;g]g7)7g
[ecPCHC1e#O9TU?d/G@=8JMSbbZAK#4^I2FTH7\[W3[d+Zc5ZJI/--c.[HB.YA?b
H^Gf)^MP7&DKLd<-?@CADO0[,cAX110.ZQV@L-U)6(,[G&]Z69bL4V1+ZS^DfVgI
VWe_Q?MR6aHW4OW5fS#H,@M-Ae,>@ecNRAZ\[^Vd]@SCKO2L&SZGF\^X]54Z]I^Z
>@7W@<0Ee5,P2<9V^HE+T)=a^.9LJ@e<C+TBXVc]S(288?.>JF1a/Pg3,2IYffS6
542?Xg0M(9Z20V0),88#b&&R#c15cQXLTdfaNY<Q/<MFbMg#[I3:^f425LY2QaL:
ZL4,X3,-UG^-&:9F<KE(DQRc5SdQ\GKZ1V.EC,QDgB:NU:BYXbU3\/Nf7J&D6eH9
P[CIT<O0.bN96[LTRV06/Pbb0Y1I&U#.:Xe;S?Q6aSA?C-4^>D:fIO&GNGI4T7F1
+6W[Xb;\S?W28F[e\gcY;T,L/&bCc3CX52H=B5_:#OAFN]EEH_)WA)4]KVR9/d=K
g;L0E(E(_/NOOgOd)K3L(GS0(25dE_]GKaD/[c^)JI6N>a=L0=@3?F>>dH:BFEI_
7e3HVaXZ.FFQS(:cP]>MI;DI;/RYYe1S9C\ReA,b[9He^+K]R(D_1V_PO^3g[eN7
SCb/^[,)[D],d1@Q:?8([5&&:KRF(5N7D5[H#>&5g)[,D?C[S<W=c2.R1&[(1,7Y
Z0M4R0&b2d/MZg)O)AS82QPGS^7HBWa)A#(N52HVL:cFTeP/gTOU+H(4WOXYfW&F
RMDf5TTE#2AF+5aB)51+dg><]P)547GB<a27f4I4K[Oge=.[;e2g]])YYLBIJXc1
1+A/C:gXS#[?]^_gPLP(_JfEJG&?A4d?D=4U5)Q3HeL?LLM8)\CV:),b#J,=IWK9
Z:bKf@H;b=289N6R@bPfT^2&a4>5O<^W7YZ.)O6Z7cTMT0JKfY##Y3M=2A>(80W.
-^edYV+F7)Ca+N:8M?ET3f;Z=+-E20OMJ&J];.D([,\gFfdW&;U7Aa<^LH<8>&)a
Y+B_6?5BdB<afG4MR,)<c[5aHb#WH[Wc+J8/85_V8Uf.XZ^;4-;[O7I^]._PaZ_6
&ME9c4:-;>bWB\)aO,D/=#NbUIUV>X9;N_/1LRW.DGM1D3V@>Ed:2/Ma-GE+A<bQ
)CCS=[05V]d8]eB[O.L)f+]0HMJdP6Q+3-e1c+AB199W5Bc_N>80BHK@<ED;6HTb
>Y[Y,F;8@f4PN;I.A&b.K_0??3I1c0)EW3L)Z[+KC?:4cSbV_E.9]-.Z^I_58Pb]
<f:QSP/4cBF6>.3R?(KQ&8B2a9X0>R75TOPNU-<A)Q,3HSZ+>S83(85d8\];SEG(
3KZ)c&2M(4QE\;a5Kb0V,QQ(dD>;&cXKJ/aGG6^Z;>TLX6?56e1/aRd_GHCWeN.<
]:;-&.#eV&5bZ11=M4#-B7HL.Tc[YgKD)JK79<U8dfHcfT8g/e(/?#ISQX/(e]]T
C^Gc8/?dWC&U+<5Kd]H<f65I>)IN)7=RB2(:cREZ?.gPM1=^ZR<:Q8\M/>Z;fP?C
-B7CJ;J4?TP133IZAcR/3::c_(2\5#:C;E\03.DJg&DG-a2B/:W7YR;&EQ/,7dAY
0>Afg2U#Qa&&OWB<YN5:-g_?3F380H-;G\/1[gN6,FT-U5f3DMY?gO0=UO6(I_(T
H=T32.A>6_0BPO<&?]b+^WHOT]FKVdQF1P,M=^GP?B2\JgA\bMaCRgZ^>H;#BP4^
=^-SYX)/H]<J;;aa<9SY8&]:I:8\??gG^<db3X.6XBg.4Z[=Tf#f.N5fbZ.FU88)
&NJ4a^T4]3(B3:B;dW-f5/K@MM:g:Y3^7MK;+UI0WS9?gK5<JMQO29<9,NSV.L67
0&aa8^/RG0;-?O,X=09(5&=ZZ\SO(QDW_:>7VN(6/=L[QZF5T>M>]A>D3&,&M@0>
>fNbfT(VMRCN/F2TZ@F,1HU(KJ_;Q^MT0BJ:AHUI,@WJU8/RZ.\JfF^P=@B\eB-#
V^Y&H-CXT+8WI7W_O=BY<Z2,Mc15JIL&bTDT:#0O]TDKR#dKH.0E^Na^Fg\R(I9a
=c)_=4RI=DO[E&=Tf;JOaY5Q.K;(4bZ8A:fG^2H)_5a?R>R#SMX[3dM#@=FO4@d?
a1<Q//M&CR-Q>YE_[#]eM,0L^]G)CEVLDX<,C;6K7Gg>0RPD9G;VCZ?-0;P,Z3b)
9BfJ/PId6=b+3f>&^#]103cWMA6=TR8fb_86/aW&>U8-G;RR4\Z\OYS\6&JYg)@6
YNKJY5<4f-,6SIg>4DQZ/W5bc#_b]X#O\If(Q8;^HET,M8<[be_)9+:g;fBafWWN
E/-M,KL1[U+>3PW<LV,8g^<E>fPbEZX<>.=#P>ODOPEWAC)fcOdY.?2];)BaK0X4
NEM/fI?_28Ec?6aDS?2,)UKVAXDTXQ@DaBVb>;V;D34]N47eDD5M6038g9BKN:X;
bQ8TKgT8\)4_D1:9^O4Y:QQ>+gF)V]\KO_>SN4,ZKQX:-G8X13WY.W,B);)Aeg>5
M<Ng24U)?&0+CP&48O9G8&(1B<c#4.3PHQ[fU2-Y7?[HA[fIK/48B=Ig4aKA8gKE
A_^>@Ze&Q26BFb6@f84:+7f6SgK4RVJ/013TGQQ2AY>(S/:VMS>3a&AE+7.6[QP>
1&XI6aaCJ(EQRP5:V8Hg1&]#2//Q3eR4AceWQBK5?U+.KBEQ#S0__R@]=F(]0/S[
9V23;6(]FN3S[QC9OR;WOfTVBZ6UKT0^US@XZ>N@PU9Y?E&0?;UT@J.38Q&>[3UN
<+IAf+LaK2B<4aM?II.g,X]?Q]bUg;b4]e\P)8L=UaE-2MN\W>c6B@Od4d/3]3EB
-)XKW?YLLScJ18?6N)LMR=[\I#[<1(/+/+54BR_Ge+U7:1d5+XLQ#U<QL)/FHK)6
B#/W(HXD66U(<ZXF=G(bN[IN6\CH.cf_IQ#@R/(U6429V[,J]]-5]Ug\:b:?A\32
9f[Ne9T;aCbEP;L_BHW_B5G3f^Ag/f5T)dJS)d5[C<dO,D#0LIaP#)].WVA?UBAg
cM-dcNN<J+S6:T88P07S#_CY3EBDeLZ_<[:TO;9T@:T=GW2#(;P/=62SZKYV@e,#
gc1GNc>KP#b][IcV.9e35P0M+_05(63.1gV)L;aG?UDg1N)_(E@>;?MfbL+.5Qa]
F<24ZHf<Nb2BW8]4R0.UK^[e]QUVPU2fLN^RZK1E/XG:E0a1_[B46AFg.4\^W9S#
Sc1e\#5c>J81)e79H[>A[&Hf[QSF)5)BN4^N3YcRf#DUcUDR9/e(SI>-=<b@Vg;d
UaeJ=(+D)Y+?KV]?@#^70<G4EV:+]4+?I5V/Y7Q4]WbdDW.;71CJ@e88OfQa0cWC
L=,gAP:82+CQBLcPT4?LeF^&R];;3G17X\gg:f>]XBdX2H77<Uf.UD;?Q,CKc&65
f/bB,RUd60_eU4\M4V5^g1@P7LV=0J_TDJfNQKJde?+W[,dF.5Z^+LXVCb9eF83H
(Z0>Qg>,GQI0T[:g2NB+/(-=0YL<#g/3gK=9?Q-/R;[;4ZQ,0&.a].4&],=OW3F:
9cg+_d>H(e3g(TIG,5eLLP=;:LSUe+W#/8>8]ZegX^,QQ6XC0M>Q6^HE,=,P:@dN
4>VRDCY>@Z=@3)XH7=3)O<)<[Xa^33?;P/P61N+;AHOf[<1UcG;^O,SAWV<K86Ee
U?9J.9AEXZ&eBZM[K?6=KE>YaI,WTH[4;,+>eYUA^dOB^1@_Y,=)IVE)gHHV,Nb/
8dX^FXFf6HFSOT0SPK.K.GH<\cQI^3QY/D)#G<HDbKQa]5c,L.Q\a#O&#>273f<+
5]PK>+_W5(B#>Q9^UXeMVV\<P@-OJ[A/6Q:([PR^@QT770?_)>;L^(>D4D@bF\2R
(YB)e/WeC.)YOEUZN=/BJV5_GRX;[\:A3=9[MI+/3@bM7-RSQB/<b,bS6YRHLW.P
DEP7>=U.=>#\8-DC@#,Me<V729U=a;<8YMGK9@(H>\8RYe,;D5.?Aa^OPCd>31YY
GRMRP+_J^a6#Z1W10TG_(L2#7ZCZd21Df<,[bbYSYb90cZZTMd[VVg<1FDQ27]1U
\D[WZfa9VXS(>T4RCa+9@2FM>0V-&O[Y:YGT3=3_L;a>:5M&5J=?.[\N(VW>GdY(
46fgb600>DY8.L@^eH2a9C/@EAJ?W#<XL]/fT[cL&RS(RTTFY#c9Da?f.L=KS_Of
@43b/=OHS[eI2U/4V_+>2YR+(52:B1O(dHAG4XFP&aTd2D51&(.G]F32@K1Bb&==
<H]++L8EWO0_:3d4IfX@I-#3P5Z1N?\#QTd0DSY2c9+;Vc<bB0MFfGM@X1<W#-<,
_TKe<A\#=\=\EX\-.#T-B[b(C&UeMI&).J_gC8FZga20S7\5)NEI=JR,]+PDE2;e
M.aXPJ6_&H#O5RT..U728(U+YX_W;19NVZSb]U1^\G\aMJOR>aVMgPX]Fa;dVX[+
_=DLK;C)^0WQKG^f:OU(Pf#UJ]ag]^(EU?E4a[g-b:/6Q+><DW9#83UDA.#?;RB_
;J-VD4[a2M>-CWGWUY]GdD+&/B[_LOV9H;SX-2<LdFW?46W2:J\-[G]S.L2(+9A2
X)VQ(0A(69aG\XI[?)LT8I?D@+EK7af)@@K8KDGB27MCTFD.Y,,HAOg,0L+MJ.>c
4D(-XT3Ne_7>fNe/D4[DW4[?HW-AgUMHZ:HPW]eX.13IG(-RDZ.WG84WGZ]SeR3C
P7TO<gOPGLA3<T83&N[O4Z#;W&ZG^@A&-O_Q)./HNd565/eATa8A@25WR#?\2SKf
)25^W5ZBL&6=0,>H[Be-c3WLfZAI<S<@F\a9D\Wc\F8OZ3PES[,c[9V#8:L1/?:S
/U^gRIP\ag-]GM(eAHEU[,V@MR6Y2OM)+7/PXO\caS#NY5KRbO=9VJa[SDa027aB
SSe.MWFXAD,BENN13Q(\OAJM:3BKJ)K^9&cGDIQ4\#;=b@^+E<6LH12H<-XHKf8H
E+G[,V0XN2?MPcdZS2dU?/@)PLQD.T(e2:;GFab_ZT<SN6R#):^FgE,G</TH;W,1
9@_@bd;/RQ(>FH^46:NI(S_C0H(UQY(W<b(3PI.P0dLP:@A]M+DOPQBb#LS8]g#;
cL-Z7R);FbK#&T1J:@#g9acgF@=ULLK<Qgg6cXWQLCC607^>I_\0?@d[A/dgGb2=
BC1DB6F.6;Z]G:Q7gW)d0fKN9#H?:f@2U&Je069D;a<Ug9AR.^R?D[-P8?Y(EIA-
XO-?8IBXE_N@?^gA/_\T95dM\5gUS=&UB<P;+G&AHPEO@7ALYa6I2E1M^[@8/J#=
d[HXgGW(IN65-__QB;NeB)/e4@9MQRc&7VSXecFV/E_&g#@XgfTgM5NO1Q[b;EI.
3_D4>B:X#@cKRJSd#:Y<VU[g<?&3O#6+NTDCS:B)Y,:Y<VV&]\(#H#E_N/,XMZg;
[E::D#@>\dYcL@32)6FO3F+13>.e6\A0:e3K\RE_TW]7LRC,SG&59;[H\bbTF21]
7f(\^Y^U&:\7?16dFWGEVaRHLdRaIfCNPcFfV)c5?OQ1K+8dWbW[U&-^2=#?bW6@
Q:2Z+8_D1f<U.Y18B=.DWTRWaVS9a9&3(/BVJSY>\G)e][9O(RV(Q:UGR/Q_8;18
Wf^W5U<.#R#)ZgHb=4R.<TKGBR7^#L3A#O-+=7d.<NH=&0E-)d.E]0K[M<AK0cAS
U8?N++cZ6T9V06g_.cKK)<[UMY],.-LIg?0T46,B]d-UE6-OV9TQ@FB.5bT/MMF0
^<e5.B1\<?Y1_K?MdY2C:a[(I^S:H0/?@B96dK+-2gJNVePH&WA2J-cOga<&[[KC
UV]>/PHaSLa0K(9@DAE=H36JfBSPJ4]3]<I(<[/ZHPGSb+(2OZLQ#:U_A-Kc8B?R
A]13J2F@J,]Y>U6-00B@bf;0SM,CH)4;RE^,D05IO/@c+62NO_Eb\e#F]4/:I_JZ
ME;WX3)S8-51X2/^8WP[,\G:?fF+CP?@baIC2[dEf<c2D4WB/V6L,/Re\:#3g_f\
[X11Q3\W8K3P\MQ:VD:/8?AAV/>D(<:ZX;FW]>ZBVc[#/g7X67:-T8)0GZHScY6/
X8N66_]QPHDULOb_ECYCE)>3C/O#2.\9:_)T:4_5)TQ264\F1[O2d@<Y-L@W2aLL
2/?Ee6cM,=YZ1_>Sd40CGbJa>4@\46F[Cd;F;R:GPNN6;QINGcK2O.FEX5UKgP@7
NF680[CLCM?8L1EP(d-=W(D;bUA>X0)YS->d5HLRD[/4,/fgf/eBBefF<?TGRAe7
>4LJZ3eGO^73FDXb9A8g)e[8U\38,bUd[?c?f>^)EK3/W,LD#E>7KOI;OYCP>D&N
+/W=8(e8\]H/5?>,ZcAEE/5&??Y?JP>N#dWB_PH4c],X3CZ\BJT@fAQU1])R=FRZ
YT&>].>Y4.?5&cB;D;..<FDEHdERTaC&R=?a(<d-R:Uf+HW]VP.:/0PZGeN5a1DG
METb)X?7)(2a.A7d4;0QLZDO9e^_Pa5f\Y\4U1,;F0Y6^AGY(V1G<c?b6g8(@0QJ
\_]2#ePHaVc_Y.#L]EV.P.Z7KK\0):@]2VJNScc3.Y>^Zd;cR=I^ADCYc03b/c59
AJcVCIfGV8COGMe0+a;f40J@Ja8,.&E;@)T)>?)N[f.6I7<1A:R@4KWQec+/O[BO
R=[_R[NQ,/1G&&B91^+=I@Nf9L<KLNIPZV.07c59=cAG.>@4U&KBfOAaCCXLbWD1
ASeA+/g#JHOOG@YRSER7G41GMF3:0(F/QaZ[Gf[K)<TNB00@JYEPQ:IA86?]:c>_
WMB30VK@NC01f:RbKXV\KSHYP:X.#Af2XQ]DY2+A-F(NN7W#NWH]dR)+]>/]G99f
gf54Fd.N_4d+3.[N28#M@Q6HH+edS/6Q1)]3N-E1H3\R7NaNJYLe^ZK0[Z3-8OO.
-adD/&MM&9DfADPcSL?<.F;^H.6HN<&DP4\5[_1IOAHR)YO[5SgUG]26K97.T,<Z
6c2R1AIR:f=CD9_H+KPTX)0.Y0NW];K&51I<CA?OP^(&#C6^K^6TH6V8dcM]b8[@
Q812\,&LI?fUa&VL3#e,3V]WeD(bdFReLf8[:\Pc3EdH6RBUC8GMZZWLT?FZ)0E_
<ZR-]?#\#Q)d/Y6\LM05d&;Y^dQI1CY;6^+,JI[3F3dNA)<g\B@.Y[#5@cA;ObO#
g@:\0>:;a@7W79(YQdgbL^D9C9gCZG[V0_b4D]P7O+84g<YJ@e2@a7K<7_a)I\QV
XQS//c6W:KCT_]TRDB[IXcR]<ZSE3DRb3fP);JD57/e.^WgH(/Hc2X,;1+U0+MP@
.gZ?VTU?GJNRbB?&0^f:LMOAI.YRJ+SL<E>Q#481/dI1)>K4CW0=+VU>PRg_b]P[
9/#aI7[.[0VAV856cdYHWLPfE3;HaDJ=8U3&M+BL7YE>1O7g,2Zgd_#UMYCAJ[^[
YfXA@BNH\S;S._&4b^<aNfGe\C8\(bBZLb#-BGQ@g5H]W26\DKS<=F-:>#\NTCL8
46-^S/#RCMDd+a?e990KD<XE;4-@fNYWJ\?L&R4BKL[I/QGAH2=,HS[+(L\@PU9V
C-g0)(+,f0EWD6c1Q3G9ML/6[82&FbGVQb/#0K;&B[7SW7RBA16ULZ&VC_DGB7XP
=QIGS+\A[YUg)Y+N.:U/(K=I:B,XKI@aVKXU/UNg1)R1bGDXPSTG\8T99R3UENW<
:N4(<Y;Z\d1,=HT1=,W#d.2-7H,.NT>0HK2J,N()Q<Q_d=dCYB2DS^L>9f8?gFc2
3\Pga=^Je3gW+RdES)BT:.g4VM0(77eXR+@?BQH@_9[V1((J^N8S/=SCI8A0/a4=
767WXU:eOXFV#XG/?;UT]5De[/,OM&C?B//)WD?PRJ=<^dMVURF7<Ea?M@6[=/18
J\>YgZ0R(V.Xc2dOZ3(MPU\)CM>B&Y6I+6DO1ICcFFX+e^^G(N@(B5?<KCI8F[Y=
;gAAb8VcY9eFXdMGB#]@=6<^^Xe(KY(0f(4U2;=_E.VN>ZOF>g,Y7eLX:PRQTR@b
6[<eAM+CaG]M5K@40H7bCU^FJ(,0\Q7bLbP_0AeN+3Sc/):#NcZeLMXJAM..9(<M
\JF_B_+\;G#G,<,G6K0B1?..bX/K/CE[d+EX+8J<6H(>2P7[9KKNbU/f[UTAP\>I
9_MBBR:YVg^43<6),I_)Q>PE7Q8[;<aTHT,g4S&_2O[<.9N&QW[<d#<@I4a2C4VS
2b2@?I;PcW@17>TE<R,dH^T1RfWMTLT0>7:K+FVgG[DLV<:f.LUbUKL.N5].GZ)g
\5PI+;]I=fL>VI/VbBQ&,W[EO8YZZ2Y6f;gNF+&-9V=HfBaJ;fde,g.-+fV:9GXV
3Y11ZJ16^,#T(\;M+V#Jc-CK1O;7aaMH_@+]9BO-F>dKQ#^;BOFIa=YXHP,,8Ja.
CE75G(7a#V\+C-7L4=B@J,#]_]/,ZccKMOVEJ7--P(:;\?e:H#W\\.e1TM:P=?U7
1=H7TGT:.<S)O&YV,d(,\>(;2+0^RI81/6c4:M1c9AJaB<1NN^8-F:L+F=DT7&]\
8eUOT.4CCO6Ce[TZ?)\(/.g9Pc.fRb2:Hc_a0dIQ]0-WJA@EDZAIaMSf;g-?K2:g
WS?/:6PC?g-+aO=YN(8DdXV<HW/:KVNNd:W#4:Y04f4RWP8AJS<b5c,Idc?0e82?
O3.D_9GG0:I6XRCODZ([c=XXb-Z?(T,cL2Ra+F<RT<@1<&Q.0b<?gYQJ9gH0M67E
SNIQfRLZP,X+JOcMRVc3FN>GL>.AZW_B.0N&]?9U6JdN=2Xd<c21IIY[8L-cf)G2
84L\DVLX\a4b9/7JY\]<9@#;DA==5CZ-KGMQH^GX,@Eb)\9I\E:DY/,Y>;(5:c0d
<?a]ZZe0D2]8Z-;/OSD.)VcJ@=a9AS&(63+YYYDER9b9Rd9UXb1QUDH1KZW^EEc>
Y>3=,A-9,KB9e^:W]UM>Y/Me-6R<:S[b>=?_#OVBgO/XML4FOOK\2AfHU_1g3JTW
/49[FYPKb:W?G.R;f.9-X/KN2XPT/0REEC=[5U,Z7eBbgg:Vb2SU)@0V?RZ)6gMJ
P#I+a0<MW#<4YQ)eE>_9R^,.UXBfPL;]G4c^>YWGPJI\#C8DE06HM/4D4-8OVZdM
EJ/=0gXYW,1D/),9E9_@EPE91W=-Z);]\c]Q+-@1NMY8_K[SQJNcROKNE4&&[.eW
D;2CXV6E314:Cc5V9AJf;=c_AfE=7QFGN>LcDdWF_OcP,MeX:g=DZg<Y<?A)G^gI
=&gF+.KG^_B^=C(S0)LN,_=4G[3H;4#:&YCK9fNS#YUN=IG?(T[:K-EAHM#^S_gd
4&W6OCN/>##ab,Y#QV?0.A)>a.HDP+&&:XH.=^J+]Q1\>SA:Q^L>-BK(W^.WdK\;
1@2KB0XE7&IP7YCHWFI15UKgIYJC?8=.eFFH98]@3+,9H7F4_c\[C]+G[1+9e^(6
9c;,6V#68>cGaUR=[QFaOX;O,>F+5^(3,[=:2Y&c[YJMQX8K9]W6K:ZQ?X2-CAb?
P=7&=GU;[?c>I;+DEf^ECS3?gDMD8:]\OPLA&-RY?5I/+03O0FF<6Od7Y7<3Ldc2
G1C]_=2:(J&4I;(2e.K/dXIG<]>_R[dK=_@Z,BAcQ9USX#&.JFF<.G8&97O=7HGI
2g)<-=J&QNHS)+7?^cA>]VFQ\+G)YBa=NDWe6S3\0XbdfLTG.CA7M0\&V;aU]3-^
]84A[\FZN4:HcO7L3ZRG8fB0/#NYRR?L1S@]g[#>MQ)e.JIF#-A(__5;H)_eRRO/
)c9@0OGL]:F+)KO4-S21?M3<,e_Y@(0)#@&/478E]M8QAX:,1PGP;??OWZ\=LgS<
NFXX<Yg5^CcMJe/34&\LR90Z=[ZZ&8/5<<9S3/57J[c)c>W<YMF^X<3_05.ENgGX
5<eO-LI-O\Hc[P.NAIUaG=OXS@+.]gSMLKec/?<[W&\7G&8dAc\eA)7N7:(L#CN3
O-H,JE4E)8eRN;1#.J#R1/Za;MXFV<RWD4SJfa?aBd-e/+^OYc[((IdEJa>VR=\M
]E6-5<D#S-5Ce:T:&)[<H1PR;D\[=a(9\X<1(J5>?Ae1Z?O/&(DJ:<7?3MFCG#4;
UF+cH&(DYY-4FO>M)0=60\5?&BED2IS:R,,O7HS7DUBc<SXH1OWN#=ZC-WRRV935
5aS/E/I,?LH7LJCL6M^.IVJgKd&ED-0Pe#c2<a@Y[B:(QI>G-L+H=@=O+>@b)-AG
&]9EGC@QQ9J,U\61XHM.,L.E]gRE:HK\O<6O[ZDO4ZJJ[2RDW#F12b04,JES/N)K
@[DM38F[JNaS:>]LU;=G#^aD7cXZ0R<3]]2L=.[#4<41?D2AL]W;BWNgGVdV0<SX
,G32b;693\S+]dd;<,/<P/E5#_#G8X#Q-9/3752N@EOCBIO#7[7C_H3(0gOE0@bF
#P9d?[YH9EHYY9E/DA-2T59GQF_aBY2XbP_EN9W#W0,L^b0E0ZeS[>]J_YRAYYCS
ZbdQg2g20e@7=Kg:X536f^Tg(&H9-ZOEF+e@c9[R,cU068^[gYcGNEgS6@GETBaP
P.\aC=e-ZZ&J=>:]e5J,Tg(83b3^B<Z.K_b)^^56TRVOMGWU^2F4^dbVa56=-GXO
M&^IFPV6F]M_?+P@&S=ZW?>a:KG5BgE9B(39LSZaEe8KW5Qce/&,JT?^DYX(<O20
N.0[DN&4N5-XD\?D/K.gXa/M90^OV/_4HH=-/R:PY#T/dCC)6P>NLcLdF?J^c&5.
O2MAPe1Y4^3GeF\.I,Ug]G&@fA<41dGFBW>-53a6A(ICR5.T)1F7FROTZR]=79DV
)9=fbDS;57X#AAZM7@FCRLOeS4OS(NAK2F:7<([b)PX>ZHE:4G#XbUCS89X69XT9
RNb)N2Ne;(L=bXdNTZOH;eb<FW<=F9/PX?@UP,#,K5SP,UGB1FPd)\(gT)1[Na>5
_3[;eHJK=N943OB3FYE,2;g8^Md?3+<OcSb+R82Jaa#I\2_E73^48I,<Ab?3E=_<
/^/.51ZN7_\6FD5Y9YbMPSMY=([&BZe+]+VGO.=7E?UB-,c_@EdS?gVD<OO&=/=5
/TBS60d2?[e\2T?O>S)<XWN?4@9+c)If[-)QHL\aK/8\ORNV;I=N:;]:OKC<&deX
<]e=A3P5R41@50=\3;dE##AcY-<_TZJ5VHUCC1IHX#b6JNUaONDd([=KfD4PbTIe
=7BBC4c4D8e2<)___/?,A08\(_)J8^S,6=D>U=SY)2SJ.d.TX40X/g+97=TYB+V(
)+[)X6J:RgTK<N=^YC#K;eUR_E#[7L^XC)NBDV85AdK2_3ff<RWL?O@Bfe7eS8_g
8Z5;?g?G.ReIH)UGQ;BI1^8JQ,TgU&1S,)I0F2+&>WOYb:g3Z6cL+ff<M?QRgSLf
P&Pf-F7Q-TfE9NJ/#D6JG\g?DU&6><YO<fLG56,:I.2@>H.D1KWf_:0,F:2KAD^J
g#=GVQ8)S?L32Z?S96\Kb37W:cGg_BG]D:GK(BCK+:).GKIQ4dX11gfMT?OHcOW+
-bg6&1SW:dI3_)FO2gS5CgbM+D5LWN),^5YF-3aH;5S8FMBWDQ\Lf/Ef;Q?EadRJ
-C:4/4G(X:,\H1fRO9EECb<G^Y]Ybd5bP1EA1]f9@]&(?b#0+>]V5ba[8M-CXPf?
WY/;Tf7W^A=(W4TeGIg1>1_@N9>[WRG?/6/.P>0XGFNG2?WL,=:T^P:&SaDIC1AA
R6NX>2[eFPD_L-NCL]OG9SU(94GE&014A6#O:E@d_7c_VBQSbK#QfeM]c7QdX3FW
K26ITTPF7\0=+P(J:#+#Xd+#ca[M1QL=Q2^B/(0\]-G?A3U9KK4)G2,G(3R?>&X)
B,Y0T&Ge[VM@;]:M[,,b=f=HP.<N.O-d-c&4DC<MH1V)T[\GF)3UVQ=V9bCN+AAJ
P0QSBFC@-E6U0?H]E.:</^UI4bE)BMf7Y.@>\bM].2dWZWRGU1gOeLO@-cIE:LcQ
#1BPNZfSP4I9#_6dKCN?+4[>6CK,>L#N#>VW,S5:ZRfE/&L2S]V_1?[FeT;[T5I/
&)3G#R]CONbgBO@YP8]Od^?DS^PXMeYF\fRQ:Dfg;MIVZI)B(Q)+B[<]0HE(NZ(d
U.P?2Xd2VRUR;@O28JD^SI&4,1&[TBA8cRC2eJC15JUM,#T;=(KMKZ3RLH.(MYP.
P6^-I1\Nb-<68#FN8<(T(d81Y)9OeBb:&QK<,dg?\94EJ[)C3bS@UWBRYL,1.N_E
GIH>OP7[1^)#QU+@W9gQ6;IAVX5bD14N0:WOV+RU?<g2S\\gGPbd^F^&,8f3gH8(
aL[bU/86LG94?XOPge\LHGE()3_KKRIEg97/<PULHJBf-e89)fRbB7+4WL_;Bd^/
[gS:H9aOD,,M>PM9b@X,J>d^=FJI^QKP4b0+5C@@:FW+M24D;^,1.gb&MIb@SMM#
NbV.22eb:(e.(D:(VB2U)I2U&FBa5\4Cd:=d+IGT\5Y:\<1.\]^S#Y7ggL)GPb0(
4Vf[P)Ie2_CGEXdE=3(66IU,<gX36])=fX)@7)@8_=VB7,aWCY](P^Ja(X)FKB:a
)e@]-;aTLNQKY//F]:5,1059&(N?\P2+7BUF(XVEb8AM+76..5WUN1_g;>He./)J
Y4BOg6I3L--(\C##.ZA;b>S8:,44cBZ[Y=ZHdP4Ngb@4]IVLU;,QG/?b_-HQ@f@W
e:M5Re^+L)C3-8VCdJ37]A)aQ?:ED,cH?3b?EEb^,CcMEV5:;c,2;Z9J(6O3aGCV
4_,9:O,Wa>1\Pa]f>0TN_+;U^0Sf5(J_L/gI58_>JEDH.BS1I-B#JcNRS<J1b;,R
N[[L<HSSe^DMSPae?c->]E_7.&O,be#YONcLc)+1U<1[2aEO-T3Z5)X#V@82=?_g
HgW2D3E1BD_d_.+_1)I68_.+ePf\ABNGbfLY0>B+:aGO#BLDD(.NfD:Qf2HTW->L
GR-eAL^,82C<3)3PZRJ>7V<Z5=@(-5D.=&#cGD,F>[;]G--B(^)\5Q?BDHdR3d?g
W5(^[L?0\d3[)9VNF[L<_+G495bRP/((_7&C00\=6g-]IIZ<dW]YTK8E.aYaVRN,
8YL^:AE2Zg8Q@7[Se-OB^@ZS(\(:#D3>ASe&gL@a6R?fC8&PIPcD2&3]cBXZ>#N1
J4X,_NGUd=/U=NfI,#ZM/+aG=3+VTce,c7:;dZJO[MP5SU<3ABS6?DP:KK#]eKI4
_SE<VJ54@B-<.e?c;8ORf83C6e_=+T8V9:/F[/EJKYG^dJ:=Jbb9D95@6;g?,Z:B
XH??A8Eg7g\[VUcdRSFS#@e2T(UZRM&bd+?:b@VbaRVWK-I+9(Y-72JH/NQOT@+K
E37D8F;Z-3&N4G5,Q<\;T1G&aWddG/IOTd^8(@D[55UA9)\?6P^Ve)7^LJ)>YRXe
+I=.].(CgXTGg.8227ge=.aY^)GK\3V;51W->9YQ#/OPEb;:b\NIY-CAf;P[TPTB
/]U0N,ND?5GdJf8YD_WeV:P==V2N28M:d:OFZ0gf<51L;aF:De#N.1ZJ_2I?b<Wa
F0O:F8A(67;8C[-0YUV)^I0^b:(ABgE0GJ;:26.d-1C^;O@Z#-#0GF2VNaH)a407
V/6gT1:+J+M31YbW/B:g11-g4_VD<cRDHTZb?0&?9[0FX0K,agP^eJ41.,]OJP5V
ON8Z<>LCA6f=N<2/KO@cf:^H[NV]gf1gMeX.[,fd])/H_d._YB,f\Z-9GECM+RK9
N(AH\dc>?XPgcGET^B-0[/CBD(64cX[4dO3[0HO).UG72[9)O;\O0.5#W;O@FW3^
#<O-#QR^DCbKMR9B6^,Ed)_/_VC_5Va@?G,<([33)0g&1,0++c\PE_G=(:JZ<Z4+
CLBAEZHC>4Z[T&,=WPN:Q:MaO1/-63E[J9d>?FQOEI/LLcS83cSEOO#^)8E<QO)&
A1=/Ta/?VOR0eX>VTZZW4c6H8LA3K(#67SJ-^3-GA#gGf:&BK>,W7.S?H+fCD?G;
c#ND-LWE_>>2;>D2C)dLJ2KQL?IYG=G=_fR(,;NJU+Z_6VNad-M^-g,7,U@3_,>\
]YV:I5Jce/W(c[GI8YH4Md57LZNTdAGMZG,OB#>3YU1<EJ;&\UcU2@L(0ZXUHQ(;
Sc4XMGR&PUG.fO4MN^Q:Q;Mb;E#K<@-A36b?I15B2BaLe,JP9IS/f^aLc.de\>J?
CX=J+/XKF0.cYU#[/.W3V.g8aT48GCE-<QUQL:HMIgQ3_;aYGZG.3gT9M-^;eY[g
,J:dN?;G)8]LM.d]:=_YP?a5BdA+W/f9PHQGA[aH+U1^NAe>?VW@B;AD6+7<b;[-
MRL#VC+N.eB&+eE(DW&V=ZBC#HEDS<Mbg.g=5#04)+E&>(6P.D-67eI7P\Bf@>E,
O#-RfR_f7SLB]YXT2:P>;Z>3e56eFF7-EUB#<]O(C(C\9>/L/dgYT8^@MQF1LMbC
gd7FP777?2Hf]#>U=1>^5(>4S4A(VMJTR_45GCD)cE&W1V>+B,b9RJ?UK4Vgb3Fe
QePTF<^cKC3b2a;G@_DU0S#/cb(-JSSC1]FF:GfECOFaS9UVf#(PFUB\Ha</D<0D
6Na_L9QNS6P[S@)[^,6,Q7U+ZcaSL6JZ_DZgf.IFGG\EIDU7AcL)RTP]Nb=(;O3I
=DLeV]3/&R&4gW;U;TG[)aXLKd_YI;&a?Cg3,VJBE4K<J3F>VKdIY>a.;_?3c_5)
a6R9X9NPg-82Q=75>TCEGBdTeVZ5T@g2dc/-/3T98P1+Ld,EPZS9QI6.V)64NSH4
IU=K_[=TAJX+I;_Bf8IQLL8D44_:eMI5AKMaQ6S6=,T&b,b7#)-SabS^^V,8==4T
QH[J>f>,8K96E2(++QBM4Md-MX=[g)SW^H#K[9YfgL(cP-)3C]g8GE_da/KO)J<Z
RRIG)NU_7I6(RQR8S&E@BQbAH\f)IBG,TL9Pg9WMb:JHM\HA0Z3S]1WW,.5fQT)\
=,=FD/8()]bG66(V0D1Y+a1F^4WH,#E_gHSXQ0d4Q:QL3X8-W2RP#CSY#3V2)](C
e.cRL;Bd\D@W<e2MQHbZaX\F0P[GW13V[XY;/dM)/1@YKdJPDV@dRcUL#;;)S=50
[;8;f4e8:#>]b[-@9_gMI9.aeNU-++MC&=Y;d7?I-?Ue&RA7#AeCNfHF(XI=dW3G
;8.&=EILc[_c[a1SZL0XY_[=cLS(:9VdgN;=1S@aJ6..5\B8.,eJBd/0(e?MJWGd
PAOZD(XaKJ@M=#V-_SL4AEBZg0a:W@SKg0FQ4+S:0We:]C67e+AH;Q9>5+c&MQ[G
b1->cV5:U@^RB1GRNEAf>6=P9FHJK5\<gf>>MNV4\:IacJ#8N[ETMQ?F=,TZZV9J
MG8_YbO69^&M]AH&9agS/9^0ZV=:V(b:?4N4F(MKga4HW\JTO&OKHUQd=@38L@Ca
_ELFcYb,eI7G<(7IfFVJ_gD_76<>FAP<?6&cAP]eUG>>.&O&fED1Z9AEM+JbCD_=
d);L\4GGHD=a7>c1a>b_HOG_8a^cf,HM1^;C1OO4N4HW?EDN(VbM9>[J:QI6TEO_
QU9,_fHZYL9F]TcMRTd9)V0].,&]eI+ZSWFKV-U7ef,1\GJ/]6VDPUJRcUX,T:RS
ZDS/7VJJe^BFX=@_.-bX^bEZ>O_B&_[-7-eJe4fBR:17JT&aPcMfTX_d:[&D<?C;
.QX[JH>V<KR-K(=N\AWeMHO:[f0PbXHJ-?d6H_OIfA;YE6]53:c-cY62_#H#]SW#
+@(KT^a;)<Hg7;NfCb=TK-M<(2R7P<?XSQO\<\+Yb3Q>[fICA83+9b7SRg,A<bZC
4QWH[43a<:)[E-R&e-2T\a#/[8S#C09HLdR/3Eb3UNK:ePbT/N.?OF;I2=^^&0Dd
AFSbU=>&2aa#B[C\OPL.;RR?2&OP0K=/-6Ub#-X4(DR]R98U^<S\U?IWA)3P#0Pg
4YG9:G9Q:@&\;AE<LS1E8->VG4-R]]38Dc_?DbCaDW[.&Wa@?,ZfB4e^NS#@VfY)
fQ+K1T#]RKFAc>6bAg1O?aTfS(6P]H/Pa318\K5e2U8E@QD[ZZc;QPKWc=gTdMA5
U?-:GHMUgP)I:Z<aR>53S8PC\/AXAaR,NRU+I@ID&XI;LI<6SLC/\^JPN>X<69W:
<.^6IfNJ6Cf.+[,Fg)#AXS=YSB^dOTKWIRDTW3TCLKECeGP[=??Ddf.83)?[@e-W
\?7R6Zc_LD4Z..ReQ7c^4X]E&BH_=4LbJHdZ_STg6)@d[CW[?4IM<6O\Q.>()ACZ
]9=HN(gbf&2^F2A&.911BP#?D<EW;Xc;T\^b-;cQWDcNRI;7275H:GcOa@VC(P(e
R+YcHAF@cN3F?BU=QK8e-JE(H[J]/Q1@U1dBA;8BG#&;)\M-(a.1;V50XV_Q;4Qc
-::Z\TO^L6W/L))e4<T=6dg(BCKK,-Bdc8+NTBUeE0Pb00+3]&0S;,6T?:^:NK73
90de/IggQ,De,T7FgVKXR:WcN(\V=I51Bg>?L?6(df+8aHG=?8S78;8[]KA(EIZ;
UO=M[,]?\[Q?>W(4M#9#MA8_8IO>V]5JRWU2JFK3Z)/c\#3U;(c=OC#a=9NX:^&R
(T>dTU7ALS<ID(Wa,^1JcP(UbK;ZQ9O(;U^=D,HJgUE)I(PE:86C^Z8EFCWC_23W
JX=fXPS^F+P#F=_7I],I^QO++T\6M_f([YU#WB(IK@P3EL/H/&2U&L<#D+M\F>:Q
E/??BP6>Zb(/#?=AEEX[SJI661U<>BA&\B,>=)KZ?_gC.9bO7e?ScTB9bS8TX4cA
OI<MF^#?RRbFLO5NKJb4[8)[[#b<:6ZC.O9WJX9[81dR\WDXHK6P[^dG/@H<(Bg\
6IacPWbNI(CF,@4F.=[dW[AaNTc.gFDUf&E2PAPOZX8<-_2M<T:XGeP8]aH7/GQ=
WWD6<)&;#)bTLe-Z=]T;U@VaI<G8YGI;W<JSeE(>WA3_bOH3X;2ePG.L.^6282eE
6CeAE/H8T]<NERd,NZW/0VPL0[;-FbMg54WKPeN2EN)?d8UUV^AY^I7f.YM<9O@W
FGYF5K;/KM1U>^g>PCXEfBLMDYe^VG>NUAeLL(cQ@XNb17F=FY)TgCZG?2Z3>1bM
32MCT,?[(4AEaC[>Ue@\8@ZY.8Q1<R\L\4WS-RG8FL[+-&IXA(/OMV_6FJR5>I8#
:K0W\SMS1DW<)c+,P\:A+DSN\a012[]8Of5YET=V<4;Vc43=M#8^L&A6W2F3B3IP
FdGDGU.P,/TZf>JHB#<T=JUDZHS)5,8J0V).Me-BaT:UDC(]:62QZ2g4T,bK;VT:
<]#=DC=F8Q-P1<APN9JA,,W\a[6]SJ[;?@G=\QW09AXH8;?#>./(1A&2C_(KIQT1
NJ_PJ=EK7,74DD&SST@#N1=(Z.&6I[a;Q01b]2O5)>?M;B?Z/Z0RN04gHY53XSac
Z;0d51Bb(;5ML41-5/\J(;f;URD1+=N-<[6LM\SSa[:Xa1CX/Yg&BH,UM6O/<[D^
X69?L@GBLH=:LP_SPENWgR5)[T(CNANO[.H1IA&CLKZOcA6JTW5UAM;MAOE(,ET)
L^#8WfB@E0I8gA6;#&;]+4]gRB#_3:WPNKC[Kg2ENQ8[/fQ18^6WgffD6CUHN21K
X\O0_F;+T3d<@O[VdL,VG@J\e2PT)YAP;@Q<HXG2F7ZZE?f](:G/L1R<K&1>VH6H
RGaD.?PeY7TFBDb>):P7(,4.2,@-^3/A<,Sb[A/UN/0&fBOJKcf\K]PbQBcZ,ZI)
0_V2-63,>HV<OW@WIZVdEIYT[U^C&)X0&ECL);:AO_D9))]bFfY,8c9ICKEJ+a6=
UCG;.-0LTM6ZVg[AQWfd&T6VU6<1O^T9;KH1I6\.;#B;0-dA#90AOC8S.#<9JV):
6C^&:gPOTH+cQW3R8PS5@D[^7IU:LEUfFeM67Y(f(W0E\6GM^^+c[P(8/O0e1E>^
DFWV_6;VbF2/\AdCCSCEJQ3V&K\bV^OYO.VR&B0-B@NfEZS6K_dXEK5P9;ceH3e/
-MZaN8LcBDQ10ROGEfTYP_K9Ec^YQ=F\9UCSe5^4AB?c7\,3)IL5(a?<T.Hb#I\^
CNd/;D;8.4P6[Vf#U&\Z9:?26+]0YW<XWV_9?eNfAD0;gUS8F)5AQ<TKcE)c3,NT
>+Z7CgC,TcGMBQXP:QY^,3,E6F(#\4A0e<.aLHVced?g]9\Q+[I]L55]6g:TbTE]
RDG&TX@b[+H_W@64Ag7aSUBCJ:Fb@G&W&0b1K]Z#<I@HTWC[dDS;,cN>df]W5R#8
QN=@2,8)Z@a[SF\RT.7#e_W@6T)0)]Q[cc[c.3Q/\DYA#,_4ST?eAAbC\Y.:d<C,
+NNDU6-\f-0,__[=M,E?S=O9R\.[[ZGWKd;F,gJ&6+S9Z7+A&LIg7E,,RL)NHLC3
>cg5UT^1gY.XKR:IT[?(3\D?):fU[L<P2GI>>AHOAH50+BXeV3]<O;^\ac[N,FXC
6TKFVVD[fH5)5T=N3E<ff_aHd>]^7B1cH@YX=N,<\g7>d1495YYD.FP?3G;dFc.Z
Q,2.c^G<QXN6V7(fR5A>W]Ge(L-bC?J#)S&1/#OQHW,H^ee:1HWaE6L4E@LB.K<G
7JID4>+,.Zdf@A(6]X1=170>/DB&S9A.UUgUR+4S^EW:#dVdOM<>]\egTFgAc-1B
34\Y7,/YM?c/@X+_K?9D@@K;0NT-F?fP(,@=V5W:BQDO^84H=92Z5U+ebHec\;L-
ZC.130S7.7gDP-Z=7P)VORTA#FTYcD.Z962F>UM;4NQ(9TBVD3@<SXYa&^W:+2H8
6<F7?@5e0I/M:>E9#/JgYV_H0-YB43A,XR]DX\#@/)]fe6N/UQTbQG\33bRA;5>a
@>/?:7^DCAGN&^?+[+95;Y0K>+W2e+A<9P@:&F0Uf#R&FG(R=DNYN1H9eBQfI>+b
SMVH_:V&&;)MM=&+NH#<fMgS#/Tf1DGARHH8F&0JY6F+F_1-9H-Xe9.<^.Q;GKC7
>_c]]I_N35F)C1#=fLQ&5bc)cBIN](\Ua=GVeW6EP:&6U]:\V@]<Sb&GQHL6#)V3
S_4G5/U_N7F:_J7I]&.W:9TT9ZJ,X.RDB4g_(:E.O9,>M,.RAc.g@:f63Y?\JPf&
g#LaW]8PO5F&T6NKX@T&,OA=E8eXXWMDUH[6)J_0OF_61Y>a5-J&V]F2GB-UG-+,
XeEZMg.E#=cO3@WP8H2=;X8\L)(]cM]^>TPgQY+XHSMHQAOH0O[W/N7:;R3^]dNR
GE@\aY@fWgdL>+XcJ/>cA2#+^,(<.SYQ;H\VMXLHP(GFOONNSbLH:@??>]#Tf/g/
=3H)>=U4^EB;NE60La>8\\7ZPV&]d3Ed1aXKOHaIFP98WY,5JY&P]T(e/0;FCW,L
U@F/W4/;B696)eKb3#.5f9A/2AK)O^g<:3K95#g#[@SZ3(=;:B\C)Y+T<e[GD(EC
^0/DSA:9G,gNFaTU^^7P9#aaBX(].D81S?B1H]cTBa1[.>5IA+5;g:c@@0[<a4@X
eaYIMU]c@U#0&(K_V3&CF[F,O.V.H;J.+R^&OdOgc[U1]N2+D)4;LE(,Ia7H(I-b
AGQQ=\W:a7MN+f,CUR@>IB5HG1FVK-WQ&&=L#cRfc((#BN>^K=M6@\8BOb8c<1T]
0/AY\>DE[R=+>eAN/:;cR),Y)a&R]aRb\)5FM1CH7FPF;1S83g)]:3aVe9(H-&,=
U_T(V<SWR@d;L-@Z6\?(2BUZg?ETb\V_ZY#Q]GR>FOD)D1IM.b^;\Z9GEeD)ga?=
)XP-f90./)@caDg8OO35ZP;VP+:X-0Ra8bJIM.FD/#(,a-Lf&S0I,[6c8XUZH5J4
b4FK+g<CIW[_Y#.31?\Lg(/]d/&;GBNd<7XCGV16X?gOG2_W6Yd3XCF5<+f]A6Db
Z^C5=Fb+^U,F&;+SD_.HUFC3P)gHO&g#edMC>7ZH#JNIcX9afHSG])JO^+@B#M>5
]e/;UO9dTA6Q,GOK0A/-?#8I-8Z+\3?^:HRI5?Rd5ID_;85OL#&8@8TH>/.FM(E4
Q5PKC(ZE@6M_93PG77=fW9>>S?[fTNQV+^bS5:bHXTH^LNSc-5QXZM5\:Va-H#J(
FVIC,K&=F)G4?YA]83TQf:7<GSRL/6Vf2TB/WH/DE>F?.=dEaRC/LQSZB5CT5fe[
>V7Xa7@.-[TH-D9O@S&_N21Lgb;YH&>0-[:078a+L#R,6c2@@\U5-/acV[<NHW5H
)IVJ+Wd>b>6;?Z+bfBN?E9U[6E3O_YDgS0YfV1dCE.?XN&R),B.9A6^bJV2fBc>G
G&2BMg71c?DMHV3[YO\Kc[cY4&4eC)PQTfRE9;^]P4S@1J3E5_57DI/4,JTXYKE_
VQ5DJ\;X]O7LeM9(CFL50[&_+4(49P?+AF.CB/OYZH+e-7a1KK,D+g\Q?CA.T=>F
H5LXa8L39;JE0XF+WM?cM_ec[.39F><V6]W5eIV^a3(4[0N+PROWb&:T^<<?Z<P[
XD]LZVS]6R7E0ZDE,^U1c/R[A74133Z\.eQO/)0Fe/?PP.R8;+YD[(9Bg6[11]ZI
IQ=:G&e)T5FN)1MQ.=2-dQVAKCP-(I#d0=d<a(g<[2[,6RDb&7O3;=#K7ac4#^J,
_98)ZE>UWfSQD>DJ?V(8=.#@H@-fB3U\G-/-0VU)H09NDPW491SH6XN=^)f3?3#\
ee\Y:<\_aZ,VWO(Q(U^[EUQcT-K#EP^EFd8dU[^LOO1aE8JfX4^OV:K9e?2K4CEd
9[\&+V-A3O]QQ3(F8UT/<.7NW@K0DLcZ^4<JFJJPT0#cPbYTag3HF#R4fAPU=FdJ
_):Q8^=Lb@[2b69BLXVUeTK+D(\SSWIF<cJ9=5<gFP[4XU/TR.)Y,40+R4DW[RO2
3&e-)\)H+a2Q7Sd2.+6U6]29bQZWaOdY+WW0RK\-I,OcRLGGfY[egCQHD<#.Pb;O
[5^S_1P)#+1bc>._cB]H-Z;I/O@:#N_OTCbN^>4B6P#^9(M#T,AfK>b(.O&Dba6^
bcQ,e8TSPaFQQ,(d2KR.QW>QRX>TWBS_=R/fRU:^[,c=0R9SR_Kc6Gg00V_UYB.Q
7Z(Z.N-dR0>D0PX.DdgYYG,J7&;b4gBEN_S;dT4B((3+V]W4?/7CaR<5ZBQ#,77X
^ICPUcUF+K\=F1IF-1d@]2Bg,-7<6CCXEZb?a.d@X(M/fBB7ZU/N5RE6F/fAfT(9
MQ5L-QUGJHEbLbP.R3dC>[2bM17.cU#L^/O4OWc5aKBa-.aRY9d,7^ZdZW^/5c#E
]NO8+HI5gC,PPG0:91U^5Q&cZ\>-:Fb<(4Da)^Y2[#/f)M1_9F^YG135..>NcCaB
5M.-\716M1KCRLCaOc#)UEQHVF)5<Vf,3W.[T_Q@A?4&(.7#g;B6)a#4L<<AO5G,
;/UMdMeN57.,A-IDR:9gJVg6G)F276;,D?UYQWFNK;9&=1T&eebGQ#9J1M2.D87K
/dI>L.L416D1D)-S#F.B.-QB0;EPd3[e.(e_J[IO.GOY4;EFFO\.()@UQ1#g_Ja#
3+^4]ffRb\BO8D44[eB(B]^&9Qd5<F8H9V@IeQ:Z<:LT[2..>@ZdUK[W[Yb<b:7M
Cf49,ZM(G.2A-I@SC=ZJPN:KB7gWTXF&A(=@([&RFEbUd&TUe/+A]>g.OSLCebNd
[,J[KHNG4;^V)GG&Qg0M5Y]J_S]V<2YgLQ+W:-f/fX(ZUZZY@Z&&CU5J<MP+\T-J
,:FX24Z.b()V,S;f+20KA[KLU&QB-KGTKFNBGD=\7PBRKXC&K[#SZUDCf0;T3Y@K
e8fI+JX>N4H:&E.CN;Ne[Qd\Ob3DC2-5A8,_7D@:a>,=3-;P,_GTK>6=4_QXYO+C
+V-H]dS.]&g#,,#27/?PJJ9]0;6;CI-#W(eYK5P.9/YWMRdYP,O7#6#f_+)/1GAd
=J1(V,250?aVFgcf.T<?YWN3=Tc9@BS-KP?WSW?1TLUU1UMV-U7E\KBOBI/U^7#\
D0]Za=.a#=?d[JBX].f>I]XW/1SC>VCTc7I.OeZ3H,FMKZ,d7DD@__(-K.X-PQ2I
#GYU=):[^[=,G)ZUI&J+9]HA\8E7&]FF;_A]?V4FQB#>4/ZdAFJ#V_8351=)eC2]
?[&1-ca/@/F4KL3#6V,gHYc1W=c^b\T-6H.0+G4(5bH7?HP]M[3gND;1]<C5c01L
A_D,Z+1(K]?N2f==/=4[I)+ZX8-a8=]0HeOe23J+e8BUGW\.P+K5]6198&=X]LGd
,9IdWZX84<K26PF.ME5>O:b2^6a9QS\GbL:Cd/U;W0&M/UT47-HbVFf2_eCXb\0M
E:a0@6I^8+RcRB=LKGNXTIKA^88,d-PPQF,9cE?:Sb0K9B-N7NYDSBTc9-4XQ[>K
BW;Y241V80,RNd3b&EM7LbBAC<Y90:/1Se<5)X=3gb]WZ=3XA3XTIPBGE5X5A3XT
9F1VG@ce1X;7T(ZA.KOE-V33#WV<c\0Y_&2K4?:&YVPd\ae=[Y+4g5a@MB,c6JA\
NN&=@f<->FSN-PMBAgF3ZOSgV_-BZ-b\P&U>=:W[=#(W-IZC1eP;cC7gc-&CP,\A
Y#E@b[Ub2W=5)QAgZ2/KO3#4TBMFN:0<PSL:8423DZa99?79(bXH9fVL-b=Y/3Qa
7@9c-HgWUX)V2)^gPG,YJRE3aI5/6^),Q0X&HB&U\G3D<W_gfXCCD8SKX7(Q47?+
4;\EIc\E?\d:/LB^gM)9RJM[G_68adNK5.L&f3U^>,<fH^7&Gbg#,>+=890a<6T[
->&:_R(B=L_+B^36+0><GI1V:.19G,g8&Q7DQ.=L6Z-aK;7MR;eL<D(7a;I(Z1F=
M[RK1M\9\J]dM9_4A+@b(B)U/J/acN0^:X_(X+<?^C)M9=5FGQ.U+P[A[3QNBf>+
UG^H^)EXFB2.ACQNaHU3I4g]01SS>baS4Na5C5R;=dX@L8-/H3:.,cR#f5[?E\e)
V91e\YDM1e-=g5B.c#89M]RQBJ7/]TF_IK]?G[VXYJFB4V;VKU-7[QTMVUR@5Sb,
-O8.A@V3J^?TY35<.]RYa&gWO<Wc<7-4.]=cOI,UgO4H4Y;6g_K0NO(1)J44IeTM
9/HgG)V&,>;V)<6R(H3R4K=+F<@@DJYeM3f^B(PCb8+f);MA>PTO_YPOf-T:413R
^K0S2TE?7T(&YEYeS?TE_;S12KS_KBAZ-UNX<E#=>K(QFSe@(_-R:^(TTA],JV5J
_)+aN3L_22KO;8S:_=C_dEXea4MG#.d2UJU).>KV_-gKf?>YBe]21Y3:EB<2dJ;[
1fI?Q/H1RPMf>eT[L5HgDV>SF>>5<KP@d)X_LTdCdE/1==;5?b?K9BPU:2MN\18]
08U___Z>2Ka<BCZ,/9;_[3#E\WR;QgAJ.Y)K[.7,YOMBE(>QG>5g#<(F)51X@OS8
Wb#;Z_<MMf@0HDIX>]@&&ND98&=faWBaH9PS3YcFbZ9B6TeR.^C=\bA9cM,aLbRZ
]5AfUO^?3gHZ.d_eXRfUZO^gHB3MN9PJMfZef_74Kc9N=(W#3Fad\MCbc;aYZ/N4
-;/AK?Aa>b6PP-ULN/QgfT+D7;0,^@96^f+a./WG8QQc,1G=D0dG2HW1BWf)0f/d
U,7;=I\409K0>?_CWd6?P>(((W@IC@2eagS=fYb;>9\29@7)g6IFd/6Y3HLR/P7;
(8KG=Ua@DF)9N&_B1>/0W^>/NgDDge(g4;O#ZQ?.MNFS4/eT11V1DV93^;f@)\=.
Z,\_OF5=,/Ob]3gEI3W=dEA85SdI41ffJ53AK]Z<<4S<dK\>(K.-&\eQYbfJ88ef
SN<(_]BK+98</)/Zf+a=\6Q79=]=K_<[LM?^8,XAD_\QNN)6@M3M;0@?N7I7CRPb
+^>#2M8H>GATI96f-_:W.;P(Q]>geTd:,OO=/<SSPO8:^C=O@73Db7A3dfGR9b&e
UZDEI&:9DeY&X\2]3?6:.[eB+A^,_fDC(EE//8#GE+X_^U7V36C-SI_V]\]A6=+4
<\)^@\ICS](2M30&TAgFbPF)d2K-SM)?YA/5OUOUKR<784804?:G=B9LO2JW0Nge
ddY)Xgg;G,2EQ7faEaVb#MEZ)bA,?R;&6YX7\d4Z]W3MEeMXcN&GX2fLDJC,JPg4
=U30\755SKNE2@(A@T#OV6f.]7/>&?Eb&G^-P@_V45XR2,8&RbB)B.FSC;/UGZ13
)XFV<>?\]9VXBNE]0V=/I^5S.LX?)J]f]cDD&-b@;;JRF4M[)-,\H6/(^2LRBBL<
+3Q4d7T+@(<V-YdJd+OM-HDV\69/g=#c6RRFNXS7WBf2UU;67#A.3-NYPXD:6U)g
U,>VAe.CM/5e71(]TM9)LZeLUAIPQ3J&^aH?@^gCCG69PUWMV3<((c31@U@(KUXd
JI@XYO@EVC,MQ:E1BCH@#1#9VU0(+K19F+PCGB>c#,#./\)8gICJI6cZ/1MO#M,9
L?:&;?SSKJ?)M&K=27JX-C+QZAWZI\4g\@2I\<a7ZIB,TTH/MZ<2(SOCMb=V&=Ha
+ZfcVa^b[JgBRH]0QS8M5&T,YKBKA=ZL]Ob4K;N^,a(N/D&\dSS4]@?3-PFaZI/&
d8CQf+<>Vd7^.LDLNZ?5(85H6?Y-bbQeG1b^/_50CXV,eDN45>N32S94A9;&4\I(
F&VD:>L&@f(\YI267UaZ8)-X9B+8I)COT#TOR8@G7]?3,M^1F-)IC9R@=S4XO;Ze
f=g13@#4LYD:F-UY4&X=E@E4AQge.<eEDMOZ)D,gI8EdfK]L2]D4:7);e#d2G5\D
TF[=/)1/YaMH(6;&#.)YfK4;_K6D(]SE5;V7SW=8fVHI;?8JEgHf7?HN+Q<?M(g3
<TSde=7J9-@]>7UEd=]a.[7daK:S5Va<)4(+4>#aJ6fUT,Xe779af0)FJ>37#-4M
/[)9FZf]@#K4;0HH=IX8X_aMc#cL3W\#T8//),Q7SV,&GPIN<)3gc8c9QPG/+5H:
/(U5;3/<^L)OgC,I0g&J;dN,/P3#,M;CW3[KdFWgdG)JAcOYg_R13N0GJ:XEH/\&
e]N/^7cE8feaI[O\EV9D)(RL^/(:Hg:^WSg6f/N]H:5g/S9Nf,CRbdXe]dd/O=K4
]@.EFQ1H1eXBWfFS)T<)AbDQIH<W#.0Q(:3AKE+Id<f<KYF\Q&[M-Q1M5d9f318D
d;da<LP67=@WO,aF/2Ta6,Y@M3RC;,,Ia#HW?cC(>fY)71F2H)/#\>^FY+X:e(ae
ee.PM.A\H@65119N#W8eA>.EHJ[U[[FEM\N5H;1DI]2-H81-dA9@:6CW,+^cAJR5
-0K>aM9L2bDI^dg>]A;bcU0@RPZ_f/bD@[/(b\(B)+O-JM0\aIWB+gUBI>S>X1G_
Sc+\Se4^Td,WR@P^gV^^eFaE>D_P5D=dJ;F5T7_bB_2H&g13)ZXG\gW;0TS\95gb
3=36V+==e7&W#=;@,C7dP9YMP_H\Mg3HCU0I<WM=c4B@2VSGV3b0KOZ07^>TD#88
KX2W;VGeHAa.XeUBST&0:U&_@fMF3&.ZEK23#OESP]ALUBG,4)3;HS+MY=Z5.1^R
4@QSY&5d_NUJHG[.<>\\[J=5I07]-/?CL@eZSY3F+fg(g)AW5f()JDHY@.KE^]D1
0:-RQ/ZYQB=-)dIN5&@WI4KU4fAB.CcEX[a7TGAN+UQ=efBHFI<MOZ_(3PP.eK=+
AQ4X[25D?<&adf&D2<cK2ZDaL3Z?4\Q;(V^ZA)U?X[YKU6>_0=Y;0c#1;U]_V9,+
8H^@_D=_d^6>I1@SYU[F1cD+9acMXD<f],/>75JZUE1-T&4D-eRF:9Xg>JMB;]f,
A4T60E5b\BbND&.TW2TCgZLaaR8BJHN@X9.3I&(Z(EF]E-/W>FK)FaOEb^CMK][O
V-L1G\Mc((55K9;OLb[?W)PRa\-d6M.?P,9.&1G=;E@f2?L^&d;D]Q_b3R@J2@\\
JefC+@NR1=PTJM1^?W]O.eX[;391R>6WU^d(M#^P<?P.1AN#4JF-YU.N_.cCR+?#
J-5=8>A?8__V)#3=T#W@)R\(e5?eD/ZH5^.d?fBD0d>eL/1PfR-&3BE,#?:EV41S
Y1UKV99EeDE@@9D7QDIXIG7D:F;YH&FS2O\Vg^E/XX/Y)R:2@C(H&e/3B0e+AJ<S
aNMIX]-2EO9/QT5/7EH;ALF+FMa13CDYDCIf;L,LgIfIB1/,M:/\_3]3cN,EO;PY
9REJ3LUHJU,TPKe@fCU8UCZV@bWVEECPe)=bY6=0X[Hb6HTXd:1cfaPY77N&7?\7
T<6UFV&N\P]OX5EY<e9OF=(1GP1adPQ78AV:6JJ=H)IS@JR\OQ)RLc^<PO;<5ZY<
\)PdGHWW@Dca]GNX0e\97=-[L<K)5GL=FU[><(dIY](CS<=HG8T,d.;JV[cD[@9c
&g;e(6.c/Heg<8N+RA;RS\c:a3:b,(]7L#W:;aeL^b948#>I;Y9/W;4ZJY,]Rg2T
Hf+<+If[g?14MM@a31])<gJ0&L/;20E2WW+,_@XYT#X=2RK=KZ41^2gPE[;f,gMW
@IXK6XTLKHT8[a,<.=ZC?1a9O0RWE2g_?9^S9&ZH@->PGDL4AaLMSN5,5>3K/?7f
_-8dTY=[;:K_8C_8d:C<f_+U8Fc>d.1=ST&EY69DT,(DFG]?Z)@L>a#\.1><0P<&
.MF<P+PB,2<3#aF;746[FY3Z3(;=47Y#<b,c27Y2gVBgE(4E/S0<0RXMC@-G[@R.
P#@bW<C0GHW3(YaHWbLgLZY<)R=5d+e7Q>a7[KR9Xg^9ULN-9ZO5^J2ERR?B(aYP
;IgRMgQ<BeMR,2@7=Af_g.ZL;Qa+d;O:0A<]?ERGABJ55-2IKY>4D7JR\FYLQ;&,
TLO7,/E@4f@g0b#>(K&bBc:IG_eXX>#DgZC#JZ=@=V6?YfX/[=V7cL.M+c7B7LdY
ROU<[1X&NJAH+5NU(bPS&J7gWW<KUPD?)Mf4UX1N4ggU^0&QeEGJD(b,?7TY;Wa=
T9JTDeOZM6c?R<5:.ZWfa]8(E/25Nb#-S5cfNEK#ceAc:D=gBU&f15+,DE;U5;eE
#2QZ#W=M915XBGg>N8&_J/JU;SR?)?F\E]M?FXJ7dD,cCQ&1#5,M/ASDTe;VV3_g
^:D:@IX]Z;<MR#48Wf:][Mg]C+QHY0P&V3?R_3#Z-SKaKY?8;WVAZd:cf..:;54K
]ZWMfFW908>;<Wb<0=622ZFQ4)S/2e2(,.B/=DE@N]X.N#d-gDc8A@&=\[&/.>IQ
FVT:?V?S^+Z.822(V6VE9:1?<D[gO_L;N(E&)+9;,\0J-a)]eR)GQ:AZ)ZGJ>XDU
X3QS?BIZ##LT&1K,3:/gH8/@[X?3e=ggd5LF&+>S:?fI3.QZG2.T.2fV=2)fST(f
-4J0VR+\AUWHcbU9=S[T@H9Z3#WFf5/@O>97\_g4=P[SL5cJ,U,X]B[cYV0]^1\8
7O@dMD/6IV3cZP^^4T4Q9[J:HL7G#I6?22MC,UNW7PRZI6V(e.dZAdL;d]2:IHU;
0#c1N\-2VFWPgd8@\J;V:f\KY#2.7:1#5J:ecQ8H4J]5](PYO)e29ad@&G-\I>7@
JNRCZJW&0_,963_ca=SRK?VS56Y(=fMDY5ZaR^.?PeX)F]))X:A0/MbOPe&Eb@G2
#_5/dEK&1J3,R6_U,g?0,?H599R8#-c7<HJ?&Xc.=SRaT.JSE.IKF6KdBX?#C;d5
b3MfR],OEW6:(#4.1N,=F21F#\cZf:],_Z844)R[^:^B#GB29(::M=[U9?gK1>RG
J3/a&)d0FE?CTI&&4^5gH++6,XVX84Y]4A0VCA6-(M)6S^8VA7^Cd_K^V6(XED^-
)8&<[-J-S[J.PDb1?Ydb8.&XO78.KXEEF#@[94dVPWOKFDN2-_,OF:EbSTUa[<CF
STIAB_V0ZR.D#B@g01N:.6681^Ue:W090J/Hd38SS:L?fX9-;S;=6/-&XSf/F_g/
K7DCM6Ja],>J_/5cNKVENT911X#6NeS5H)CTD&M1,b,]OJVKM7R/be-OKS#]Je:U
=HW,FdO2<MD@g;[R8D0ZP6\D5,B[[L+JM\b^7;Pc#0JEJBf&S6b3c#92SOEM33D[
@EfA<-@4.7HA]a@D=Q2LT;=&9S9,TfgHBIFA@egIQWYSH,e6aV@_/d//):0[bXN/
=)44O)GEGF&SYAW1^S7&(HK]2UV=Ka<6CMV:.(C;X9cL#]B3G3Y(efBg)89XH#f1
&\_4D#P.B-e:K.18.Dd#)c/G3bSAJ_820L8g[;Z_3.X5_A.UMdS)^]\NDNbV;>Vc
ZR&9N5J2=7T8;HGN0:\PcE^>(:_69P-c3Y&\/_<,HJ879+Zg]@M40E;;YeLK(^ZW
)L+=\[/-KXPG]8L_KQ/He06O]9XT&E.HLCH)<X+<6gG:46YS_T8E<1aA,02Bg__N
\WG9daX&I(YB161&Kb2B^S-&_f=A[,9N.[+T/1-]MK:5Y:a>RIFYIT1W?@ZWa77\
9e5D]S]\T)70NB0#Ob<_SAO=gJ3H/cL]>^1+32>)KHGKK0RJ<=)CPHQ3HH.b^bD8
9_?ZFF,+M=?5A[FKCGM\@bIaS7IUV:@DY:^^De8:>Z\a#R-1NRfVT2g[+Ob]?[9_
dFRYQc<Mec8?9J[R[E.W#=HS9WdKHV/=K0V]b4B/:3?Z1c;C#KS--PS_3HEK^+/f
5=Sa-:[(.H0>g35]&,+:HZUF&c1]XId\ABR(DN9LYLWGHc=2<G/3HV2=M(3=VRbO
f<\bPJgJ/VaQ]09aZ3J:@R=I(gQ8=e7P1+TLI5U4P8/LW4DUgK:^7fP63I6TK)Ne
I6#NYP6WMACM[S5G)B/@B+3Z&/SS<gF4F8e>].++I77G>L:[>HaNGVaEOB>R[?^B
DRQd;CIa@J6MY&,PE-988b@150(/^TM<Y:6cOEc-?AE;,B<?,#IaV-BSfa<Z:9QJ
(V:5f,f=+0@28ICb0+,2?.cN&?-<\2(2e2b0(>DPU:bDQ_F6DZR?@0.IJ9&OIBTF
0,agLI3bMb(];AG7T<AVS)8CF\Db14BP2,0ZS=g6]8EF9_TPJ))I=:[]BI?)O^):
O7.gB+304bX^geDJD7eKeUcIeb=AP-6G0@U9?cHZSV\Y;V,R>,&7@R15F5+8HI[L
dH]gDa3-#a1T[=.IWOabRPO#69GfeGN_<L+TL8?<Ga+XYf8K:C;2eI@)XB6+V.eT
.TPBG+;23\#2W4]5_aZ.7f]D&,72#eWY93c8I2-9B+:7Y;OJDcAc)4]]6_T7CgO9
e06QEO>[:f\LB=/a]TWB.U4X1Z><AX0@/dL@7@=<a(>X&M=?dQ:cOXUL7HKP5?_4
8eE-E.dbF5M))J(AEgLA-d=^+8)gaI)[g4XdY1Oce<R8?CegH2&d=cRKRKPeeI_S
e.@4)C4BE<LV1bU2XX969/,7LGfAV3;NMVIN5@c=2:<E)0CWA^fL1D@F,bJ7#M.-
TC>&KE?]AYIKBC[6#()FH^N58fe5;))?(T6^d/INL[@5>?9S#?;8/#]U1E[DCKDF
bEdCGFZaU#_D^Y?OEZ?]P(#=4>5>D#@LMMX=:PT\]aYO5GbOTQ6E09,d[Lbg5Ya:
BM,FA(/NFe25<CS1aUN=:40K+(SU8eT(cTITA7#<8(f)18;^^GU@J\RDU)(]D2QD
5JG#8W1]#a#S(S[3A6VDeY6@>U(U;I6+U.QVG)g)?>K/2V=8,dQQ(\bT?:+L;-5/
1HG^4d<Hb@2V2b;LP;<^</#KM16>=E-Q3H?0<PQ,Wg:F]<a&E@\E:eA5B]>M]HMO
ST^R[_9XQB8Kf4Z+CXd:WJWD>P-[dM0]ZN?_-#TZ4R@Q,Y:;S64D<(1;>gf;c3W^
:J7PZ[b^5e&#Q(;UV[86KYe?U8@CaWH>V:7d<dM=;^1]T)7BdD)[]TLRSNNSM5B9
PW,^TVPL;B62,/P>#BM@&8eQ7dTf4_d\+G:@<^dFI07O9J4aMS]/NX@#g3QD4aOX
SI@HELI^CM)a3eT<)&HA495O@<^a6fFa&b3O^J@VZ3<N=HV5XCa[8<>[]AX;CM;9
+6AC8Yf2O/Y(gOMS-=]?AP&3V&bRD3PN-M(3,beM\IEf;@;]aS=M_>QB9Lcc2?HH
a]7A2\2.75@FE:<+a]KNT6@881A.OTgQXad.a=BT63d_5\M/)2)[(9G,fK#3AE1>
bfPgDKR>EbK>[Xf9M#XO@:4Of_L0@6Jb[98c5c7SY?R9,^Z.V<2/)c1-gdYWaY=6
>[XL\e;E<#23[SN;;\g8SEA/Z@:&[F=)5^DJS0f#D:,3#8;^<T84c+D\Wf1]9-^.
g/^;D,#ED5^&ed5&)F)))KUK;7D@2[_V3fH/^]D(6[T[6E@8dF+/a:@\GY+I9K&b
>Hdc;:NZ#H_)We:0Y64CR[5X-=>(9CNFb<6+[UgHVUPV^A;C/<CU=0=a\+&)=;Y;
b,@__;N@Q[U&069.?^]8.5fZ+]TY>]IEFTP]GfHV0f>G9K]3+(2H@R4:Fb(FBd&5
#JP96aOD5#K2G3DGCUF2K9VW<XQ27-8cZO@]JcW>77G25N+g#>JKe7]b7]QfMgGf
db-8NHQRH)<MLU_.(+_+dEA3)F<b88CU^.Da^.5PV5]4R+4ed];<#KQ@/K&WI3d>
9?.e&J_e3IVIJK<X+(:(/;=Jd:a,XC,3FJ-28YAO#-K;L)F=-Y9/N=K6c@-7YbBS
BT?_fOY2cJH6DYCHI74NRbNIRJdGA\bO9<^aQ,Q]S#1PO#]L.\PI>N:KZA#&;[Ig
bS[+2e+WF0dXN]dE3>bAYT8<\KE\K2:>>3#.;CWS4:b3NE_3G9#+6_\@2);Y2N/W
NA?=V7Qb[YHLHEW8,^gMOD]D^4[b?R((Z;Z0C@X681C9[Hd9/FT_13@8V5@2G/@I
#6W=.UZ,N3C^?WD<)T:Z]]Z4dgWc/&DLea>V-_D(65Xa9O;VHS[(AYaIZH<X\GKa
1[=a,T.,d?ZZE3/#A#L?Q.:UG:M5QO-@S03JeD4CTWP]>SI50+Z?gC@YJ&5K.3c+
KT-=e9W_R3g?/.)a?0.6VE/.IXE13/ELbJ+faUW^[+/Oc/1W;:]GV1a7-U+W10=+
2VR4<4?@BMC9S7K[P8b)eF_+[8V2a:XFWQAH&&>_9-YZ-RW/9(e#+[[(Hc^/;C+T
4PeeW(7UfY080JPaBgW6;]899OD#-6<bEHg/,O47Mf3ea^)DZUUTZ:aA^93ZLUF=
T2bI;2RKI-KW3;?ZH\0NT>8:bd/f&E7_M);F^^/[?EJX(=W-A)PdW9XY36Z#1FQ\
gN1YgK1g&,CNHd?FN@S)>B#T2&b::2&76bU5=fO38)QFfG)KC&0_U&cZ\.?R0UF,
c7:f-dEMV<M?[YL.>(6FE/Cd=@\G.)87U.3(I0X08Ng.O[KO;+^1ZNa.42b/(<L]
91VQN?gNeAO[>RRNEY5GN0653P5eN2ecWc\a?:2Ye2K^OG><M^2c?FL:?KJ\2cBE
eNB-EC+;?Ec/2aEePD1ODbA1Z)>L7(Y[fN(X:JA#;#2d#GY.<,0\F@a5B(I&CD[6
98(0,<:dXNZK\>(T/c5>W403ZCVBAQ,JWbCG>O?egH3+FOG2O]BNd<?:J2==FYF_
3A-;bJNP@&>L9&_M4PWKXEaAB5]T/F?]O<5WHVc],S5[dW.D(8&aS^abK^G^C-\X
/\31Y4M>JK@Z)a\KPeUZYXX4cO>;cL?UIGEBR]O+:893Ad^NQL+NJ]X9C50RH#=1
I]YPLcTZ.UTWSK0O^g(?\5)61WbEXJG,GX;N#IaO.c^d_Hd4:]?L=[<V>QgTH>+P
]113\dN4_E8P<<^ERN<J/=CLSN]EBdF[G5:G>4GIK_PF5b>+^V/5[0+Og=a-D8S(
A_eFfB\;Z)V<_#U(\bVN-21OMdeY1ZN)CTL;R]#)9?;8K4H[59UM[bgPP]aZdXM;
SI\SS^[;0H<9XMWY@5SQL(3WG.SY;A:?.?<8RM=#S)8N;=-#A2YJd=(E08]X:S8?
7<G;Z&N#ILg(53afUYA#Q#Lf&5_)1BZb-0-_OUNg-2A7-Na7);WO#We:>-R\5,H,
#Ub<Y2MUZdb;T8PX2)6dYW<)=ZP,?XN?2Z/_Ma3Q\9.X#3/>2&QTKTg8Z(N73f3F
<^e7>Fg]bN+NC7F4K<6^EY56E<S5IV]/UA)I2aLDUWWZI725HQ_A2M6./_BL))W+
<(4ETRK+C+9F=VEQ[;_>>G,HG+RF[7/+=f:Z25Kb3bYaW\F(I(AXQ.EKbJAWKbYN
5XFT9.U2)?&Rb0)(@D#9RdHe/\L^RTPJ\[K5&[;Gg?G>STe5L>M(VS[7#]=6XH^\
+R:WURS9)+CSTH=:OSP92>=8BZ0#Kd\\+6YHe(TZ<Rf[)7[3:(KB<^\)G?7a@=OY
]71/UY^<3f:-YT,BBd]+I4-85,aHfBY^4>-?(F44P4U:=bQO>1=B38/F7JT/)HBe
66f_63?eKW)-&Ad[c/H(J=:UHZbN:3^C>Og8\e8\+?PQE:YJ+>F2PA2+^6b8A7Hg
1A=9#7C)++Mdf2C,B(02&c67^V2gAH_^fW)>?PV>S-[1g7O;D2/\WKBO[W+=<Oaa
4B\Y/d82P\SNL6+C)[V\C,NU5,(/CA=@.^IJ19V2[\.10,R7?1cST#>QXH>Y7&E(
7MT>F=cTeS/\BR;B7_O/GL^VJD7.]ABA19c.2VEK2.?)?@_A+Ne6G@4EW^U@W;@A
^4IO#D(<ReXAX:>9TB<^:ZPZagVQ8K+f.RY^,a<VJKaS+Y\CNBAF]9bBVZB\<0JL
+\8[ZIaS>JL0M8U#W@fb3NaIW4UH6HR;EL,8KW:L.9(XW#/:GTLe60@)&479)VG&
gD[20J)DfRc=:A6->YWO1gaD4+B:e-D]SI:?=O1cT3,/CR#b#F5Z-#b_/d^&dMUS
5WPAH92d)T\2>g\S(L2CXd;-Q_J9]fTDV-,W<):Z9C<DKHeS<NC_XKKIO&eb83eB
2dBcC-ga-6=#IJfTY9_Oc<DZCe6LUbPF2@.cC])-c--X08cQP/f3Nd-1ZS[9>[,@
S9JCJ2-F,,FCDZ13\aX[.TcCRR2=UR-Q_OIJB=IY8>OUDQe[8TI/,92OFJ5fIU0K
04OGNXJA0G8@8L#^eWK+^D]?3]_A<d,M3BQf]Y@)V9Ta4F.&5W70SfZ(QO?bHd7_
-=;bA&c),Zd,dbHc(>g-ZZY;J2L5F0ZTSD9\&aI:g(?1/:faG5)3OZE2D[#\B6.b
0(.OPd_&=K^PX7O&g.QM[4cAUR7\WEUNC,CX,cGH1#UYNMAZ_WLX86d_ARPI/I(F
;,4()PI14gE=8,43U4UOc@?MOC?]cE&Y59SQ]b,>:=,C=)M;Ke6CcV&:J]-cATT5
5&]IMDS=K=CeNZKEIHJH6aQTS^\(\:]D+73GB-#HW80AW[C>\OE1g_,U2G:?^X0+
(DTB/A3O-SZ,c2WK5ZN4>FA4;6SPUGK<@0ZdV.&/_R1?;AD])f]CgOGbdb7G2Q[9
T(WSX)2g,Q/@6N3XcN\8?1=>#8(BE2]ME(@KKE8V161>S@&BJaH/1M.0c8DW6WPC
PObOO?2f3B+79f7;6Af#V66W>6O6-9?(NZ8B7^OTU1_&?cV2^A??\]AN)>Sd3\M+
(,G_8DLS0@=<F-:cU5.O6+@.(Ida>5K<W8(7TP^+[Ue3=IUQ\MM:]Wc7XCcg(c,a
a,AN?0<eda_fa&Y9@,Ve72H1X.OO4E34D\,-cEd-?=G:UB)J0=M61.>5SD:S;D?\
D/VCef<D^1+J>KUc^.PF2QA;36@78+/^fNeN,VQ5^SS22VUDC#5P@ES6(e]1VVT=
f)1PIeH7_0-?[RC@cR27Z^RRT>#S1]9J5Ib\DXA2A>Eb-03aaY@NYAA6#BMEI4aW
7gP8BYWX3+UV^.8b4\[A^N2ZH\2Q(,7W@XAT)G;N;<7YS;JVG^NA^];SE:LCdZbI
NP\dBOM(^FZbY,F=45M[K)D>Qc8AXW,MVKMD>#N_HKeXf2_(33a\W?<08ODeHfLN
:&^&VB159WfWBZ[Od9)2\M8;AII,\U9SQO9f.5#,aE-@R3P8,>Sd5Y25b0ZR.?/5
1:,8[<TaVf(PdZY<^-7G>[=X]WID?KDYL_A:D>93<G:IM.,SE_V6GHbQ0&/dZcge
MbS7Z(7L=W/C&7831R3G,2HF^A_RZK7Cc/9IOM=2X6<+OdSJ@.W8ZR^QM?G:LWGI
=/V,65//>)LeGcMVbW.+?N4<2OTO\N/,(L<;\ZR/b:V)]N3d57eeA<W_+K71-/dV
TVF,KF6I:W+V?T@<bZ2URH]&,58LM=937KHL.;ca5AQA+5b2C/cVQ)eHDf,].gJO
S9VXC?fb81b)Q<&&CAgJ>G-1J@eR\)K;0:>d512O\T3,7+FFc2]Bf)J0\9TeP2O]
T]9./C=_V4FgB_&QXTHfd>Q@FeXLf9QNO-fa/+6)NKP8M6H/]5NV->X#(8a7U9cX
7gg2;&M=QWfb[e)[dJfJV106P<[?E0^()U&/>9R94/U>3ebaS[W.OV^]GLJKM6d3
P]&K&ZXZ,=9)gC9g6D@Z=1a-;2>+A@beKZMa4+5RcL<MMAd-7<-C[9MG;6Vea_<f
ZFI7N(]X-cMda5N9/34=eY+ID,N_M1V\.Bb4=3e:>ZfVR+YY^.dCK#MJ:T4_[G8;
;XE9EW8MUb#I0BSD]U\_75gXBIAGJ3@2WXP\,^543RdDH1gO\e:Z\PVcLZM4&/e1
<@b#LYBD6PBQ@HP6@7EU^?^CT>^@9^WYVB>eNA\aX+SSD^9U>\9H1/;S&gg:^(>S
DOWeQDOZRV,44\C5.bH)GQ3O.;J4MT-[UWd\F-K4@DcWg>[;3gO,bPe4f]gI[@E\
=)KX+AEXI=]N.K_fXD,PAB8]ZceZMbPG+d^>Z=FT<HacX:\fH6fTKEI-^IQdb,g>
V,Mb:Ig&-(=@5>_/<]bf3I3OdYR;S99-d4f[3<#a]&_5eJ37\gVaWHb:f0F0=[L2
B=7WKEX58SYS]K.[PdB+][_ATQ5\d:1Y--KI.1R3>JF6(;:;X..@2F=g4=NN\>f,
X7JG^)1R^TO^UE+H-fTY&])C^)FQ8B-2a?PS;7PU>XL7#e0Zcd0\M/4WR7TQXANd
\1^.3UcO1VFg9KR4g@.f.A#GU034[LH>(ZYK?8M11b1H7SMRa(Wf/:J3CXM&J;]7
US6+_?\\&CN0[eIeUM=[V:He)WEE^^H=HHN-]U::3Ud@5-^5eJB]2gRQ&KP#eJE\
7SdWC?<c?BO7ZCWJQ63DZeB[7\G4c<g:>B3Q#U]>G&b0>QN3\L6-@HB0?1B>>1,<
YcW;2SeI<FNf<U&[-]-,]7-P>&.SG<#ae50+]9dD#92Zf,PdSgJ>5NND\<MDV#)E
UUW)^_)<KHX_[Ec1QQ=N+^Z8UJBD@dN>V/HHN#YH3KeFgNcb@VMX,5T;Z2R0G)GG
-f04D0HBBIIY@<:]^f/84,YQ&=PE:]KJeY],=@\PR/TXX.#4L+E?]f@,T_P+.OCK
X6e.E#:4>9M#.5Rga+O?]4I6A;FIaV[Q##gKF;=_g[USAJ(/IFLCXE[Md()@#UXO
Wg,U^fS_0ebBJJTECK_B^0a8-:/]6..,NI/c7;[:3??9d0E04C81g_IUY.R&T.e<
g4-b3R1H78d1JCX.>^/Z0#J?UK/08-\V,+W^.K^CdCc30/N8dScZS=eRUAe1-TEG
g/>VT[4J[\:W5GC+-LG)^88WI^Y+E17QE)8(P1ETS#aaZZU9\B+fe0XOMca@b&^F
M+?]\+PL:A7EQUK=HC\Z/I=0_OX]DQWbUD1g8/YKD3)a>\,6WM3N@g13?VS+4gYO
\2_N6a51YQRSZQ7HLG?N=S8Y_b(aSK5:VV,Ja7\+9VfSS/O^@P;aTB8a5;2]AbeK
Ag1+YAD5##Z>a:#J]4g]]f7:2e06g<Va^B(c,VHYaMc,OSf&M2RU2g;73e8O.L-,
118e5L/,aeEeYcGf7SQ(/GM&O\WbL3D)Ta>+?007=8FJa@/&40)IHZT1_e&9L[d\
3:6d10,d;c4,.;U,_R/JFD\B2?9W(VGO3C0]QA8/^)9bc4a-B739;5TZ([D,F(aZ
:[X:QA+MUadM;I>2@[XS[\<ZY>[#G6O.?7E-OEb>f]Vb_T90HD5QC=AL#;I\RcS;
>4?UTHX&LVdN3c6ISRJ<E^O0d0BVW@O?61JOP)TZBg<NV?\gg2UR#<(6b?C^;BEJ
c[PM0I]NE,T#^1^Q=g3J^a^A029FN]_X);U[YaF86&JPWK9@6a&2,F?H3^[K1Ye_
MN?^(d^-0f?WRNF+ID7Z=e:ZQJH1QKIT@?<(0d8g[#N((;Z4A=^855#:2HK6+RP:
))M@Ta@YcbfS69CF+>HW)ac8a1,Z,Y##XU/KB3:L=+\8bA_,Y1Y[RLOJdP5^Q^S(
bB2fJU.;JSW^C\aN3]8_BF7GO3Q])IeX[6]f.HCM)4dCeUfWY_S-J/Wd8AP@J@7+
Af1e(Y3&#8d]/RO[\8G,aNVgGO:B0Z,PgEJT?;9EOP58,@6#fV]670#g,1(W&W)e
(Y&5aGPK7a4E/+6,d?Q7DX((EaS=C?^@<1_aA,f>9\>-M#NNZ@bV\g\UF<>&AE^:
dY)ADg62,23+T-?c14F@:YXB2<7Kb[D9]@f>#1c/20Mg4N1c^/W=@A^01e2&N[<.
0X)_SaE&eF_e&JfYPO?b@&9_Q,a1bTD>c&XG6eARMQb&#DQUEIQ7\Z54[K4A^5/c
\]BF;M760PY8;6M^?f5fb\ab1bGC8S:H.ZaYBgQ^157CGQFBZ@fV/R:(d;-76NFF
.TGR2W3RSBK_Ve)6)\I1^dYRFTB2f]VG<^7BGcG.-fA@6.X<28Ce7e4>0:]aS^_U
;[BXa)#2Ig2_f]@C/0g6]>4G^1.@]d5=&+ZKJDN+.?bKI-]FR/[:?[e?M40cbN._
P.&-RD;Bg5-DD-LY042X.:<0;SP^K=XCG3S(E6CB;e4SUDfEMRef^G;FB;4g_d)A
3c[>[P^?S8fI]S0GZ@J(4>>-9>,#M[IKG)K\J[g1XG:,)d=9/4DKSeW=-DJQa^1L
@6[:5?W6GK60>UfgbNZNc[2bTbXB##]DZ=M-MAUF>D:EM^Ic0:EW;Uc;La;>]D3F
acIT&e9YNHEJ?XZ7c/A\&8-46M2#gNPM+5<@K(S52F&C_#P11933g51&RD07K_aH
1BL:VF(+,;WA3+(e2B.B#BT[cJb@a#\T1N^7.Wd<.dVA)b^Q,\#)DHDO/ed51Q8e
9G>1&72]gH+)(Y/;B@df..\KZA0A1^ACLaE9bdZbJZU4g<H7PA->Y5:0A@]97Z?d
/X82X8URHRd-4C:US<dfg(:QD1T_e2SA/[[=7EKDG_+?RYVXN_Y5R(N.LDT?Q+eI
8c)SK,+P6/^)&75L\D6YCKdJT0]?Q-&R5P<;>U9NJ;<Bg9_/MUDNWALIa_f]D;77
dGadNF>0MO-C#aFS_FQB/FEHDbQIM2]AOLCgD(_eKe#[4BTg7YSJ)/8Z?a9>#=VH
B96+<d,IcV?f+4WN4fQ0PbY0+b-XTQV@&#84NZ[/F1W?e2#V?0,6SC<[L9F,VEFF
,^BWA(gAJ/=&ABZVT.,\MeeaR:/8^-Y=c(R3&aNR@H[fJW^cddff(^a@DbL)KIf6
&1H6fcfWX8Qc0A<dg^ZVC.,S/Y0N\N8bMX&#7g(.FdB4Qf7Jb2f_,2AN<b<4]69c
2[C(X;VH.K/3PK-R0cM><HR2d8EX=MOcM=cfOe(YTB.=?g;;YA.(<+#]&[]^g[cA
#X6[JUI+=dC:EYBea6EFE#(PG@BG72,BN]Y:&cL=Q;XbGHHJJWQ_XOW3;&&5QPZD
LBJ6^/OF+VGTYMFb1>/<])R]0H.6ae.Wc&QG5D/0TNC\5_Gb[^IV]3.4A#,<U:Hc
=7]WKIYIf5&6VVcNJI5NJ3BRaO8)\4BAHP7c@9:H<QUSETV/_b[T&d5d)WL[C+_+
?JP4dXQZ&U+DK,65+CF_1DR31VQ&GVPQB6PLJeJb4)QDNJ68d1:@?FR-dC2;^=WZ
HU6b<D.bX#/bN-Pb^5(FEa2RT1Q)7^Q+#5b+J&7NKF05LS&>ELeME==Uf]f,Qf^#
MZ2_ULXVCEGXZ]5567Z;S^P??)R96(?3UW&R??=4ee8HU)XLI_Jf1Z-8=TNK^dg<
MfG/&JN66NQ.)1:0<HPKISX]aPEE-[HD?XgVF,SL4CU\0PUcW#@>2f>,d48TfgGM
HM+a1&L)?;+(NMGeQ6_;@+98SZ-L(:JfM]gPLXZ;10@4XB9cVf-KZMU+^YO;UMa2
@,,bSX4AUf/_B(;WfZ5LYW:,KeJ:Ka7T\79dU-T12;3f2@V-dE+0))\KbWHfbXd8
AL-G-./HIeKE5\<VB/?KdX=4AKJJ7DQ6HM[.]X[+./fI\PUe-[_[W?X<9c/EWQ)]
LO3?W?J:P&]BR2/INV=S+K6fgQZb&24;?SLN?CD5(\dK9f7M4G3D-O]=Sg9M\5aQ
ZgBDX,Y?6)>P#VQALb^dJSWW?7a.4)VCdT_ND@ag-:SF(S\b(K]7[A&UC^;J(E5;
8O^__If)d9B=\8PB;^_]2,Z/835,S1ND<bS.bQd;.5CVAd(79PgG9RT38c55DB#[
1:031<cU@.2A-ER6>]I:0SN&Q-YL]O_4;/dG+#4XRCD_D5.)UT6DU>.[8J8I7&A,
GcE34VYF8Pg=53/HB8S/GBCJKKBZ\ABOcNVXP),=Y+5B[YPZX^.TX3O4D,/0HC@U
LLCbA;Z_:PC7<[/F@fM_()&:;AGdXA3+PJc9V4F&X,[.V#eRNeP)ZGVIU[bCF34c
0<5cf2-@@dI<4a(RI4OgQK\>;\-31Y66JW3HEV<H20Fe-UfUODCKP+QV4K[Z:\UX
DO\e:R.d64HGX07I:e_FfM^2JH<P<9_g_#:EMXJ?=L>[UIB@)4aR^f_S(/abYMgL
P(c_Zd<bL\8]&E.Q5:12L)#\Z^IZ1#&3db;8H3)a\#C3])A6OP\^_R<7(G9f76[^
JE8<f92N;>Ub@A1/I3D]&L_VI?.P=^HbG)S8KMU-[:O73&\61KTOcb/GVI/T:;g^
PEaSLH:C(b:@RKC?:>[T^)G;>JXR<PcBa]:06\R66eEK1e<@FfG??^AZePU\&dM;
GFBLb:PcYSS[9Z]W]=T,@)2W=M#<Y97e22//SWGC4;]UEQ[cN/:5=<].ePeTI8<W
+.E)TE@)\P9E3?VV.L/L<b25b6G\GaSg6TULHRRK_.D5O3F7Q]T^QE8?[2O_)=Tc
F-_I:=.YSPW[L28DV5KANE[Zb,fU_0?G1)5(-/#aC/X.TS)BAEY<(-N=8VOeFO0K
b&f5EbdI)R^7?\60[(/?a.1:;^ePZ6?K+#SOA)F7,DUSN.29-fCgWF_7,X,Hf5G@
d#00G3PA_[=+-H:2A+?)[_@FNC@?UO&a>#+3-22R^dD1U#O0H#d9_;AKOQ1R(d,Q
-P<(2#H6>F8(P1X&A0I&bU:&@TE7Jdc39QZA61bVO^M(&.W8O4V&4TAEeH<&aD/C
YP8#09>_O=PW(CPe+VEH;&_3F]-eCaf4YR@=;?ESQ=6OP+-7PW=XEga4X3WJ24._
eZ8[&(27D.+[bfO5UHPTMZQ3Z-9R:F65Ac1dHR@MfX];S0Ra_WHe?d<g6HeP30#]
(H05=V[FSYFK_.52AB&FP>]eZ9_\.JPe+cD[1YUN&.)\f[IaOX.CZbE1K&-U675P
<e7&NBQ\YU97bIA@0GKJRg#R\LggbGJYL=&NFK1@@.I.LMeNX>GEI.b;,>4/.U)]
LWQZ>F4ZR_B81:1EdXE@4C^.W24+f@I^H5a<>_4>8f/d/2@.P?E5EUS;HPg8UPCW
<a(H2/gc3OX]c[C]9O_O-U+.BDCNWef>K5=a<OARefJ6+Ob=JW/bg\DIEgP],([_
6?2ZN=.>9,?@ea)B,)YV70&IC<VP6=ecONE:LW2C9]^Y,C3_PPf]NZSdeXK9YaGI
XFN?TCA2?OaHX(d&(KP97egGIQcO+gb#^]AI2OM_K0<>);TZ\9Xd1_Jd5]7QSJgH
dO&:SDF00T5#fUHAS\C4MLc^GcQFD@76\d[/^?gT7Ze.d\eHb7U7:)1,5YNY0SE4
J7,2bDJORXL0&ca@1;2L8/914S(_;YgQdE#V8XY>X55_\(7:&Q8IC69Tc596=IDe
NL8[(Ec/^fBGgZPa,/&5SB0EX\daR/dVG#C[a^GFV]fC7)KTYE3:,J@7^3#3<,&X
Ec2e08>dG.KCD>^WBfg,e-]K2WE(OccN2LfIGM5W@f-SYB=DI/VI4(.<Q[@QZZcH
4NHd.DKB54eUK4O]<@RVJAA9?WZgSa)PQ;7IVAFN/fZL@_C4CeFP2Vg7+F,/#<-(
4Y2e;VZ74SKc[]bagS@.cQ@P#=_3Vg9>EN,B6,^TNd0b_;_MOMaF8f@G=P;9CDWc
\RE0-11LK&5)&>;A8G0a[>J>#Y>fV/O<:EQOOG+TA32+PSPYZ3RLOP@g]9;85,SI
\??72GH2[E&MYF>8M)b-SGf;VJ[=R6BDT1+#7&2SY\\8&)2,f0Bb(L=ANGc(9+UL
c#&ggbN+T?=CQ2[(g:UB>PV@JII@K2/2;S=bZQ.=BL.4?LIZ?AI(S+:ZG)#3WOga
+/^C@+ec61.64LggB0eR3,<>g\GO)J11WZQ0;^I</(^9?45OcdE+Ud,?.#K:gA+W
.OG?<B,cJceWaA_GMcCU3,?dKR3f)a=<X^=:e#c1Zc.,fFW;@6)Ibg<LBaI/@RJE
77>5)I:@Y;<Y4((CXf-];J\?)J.4gag]W6J=N\H+OKO>;DgF.bS&SQ,JR=KT?H6f
7<T1NH57f63-:De43:Xa[[.T(gX:aM9[#,A>QOL_=7NR#1bF.:)?bNA.5P1MSHEB
_-eLa:[G1&<XOX=-ff@W_H+O.#L)I1;<8ceZHU:6X+]ED=a9GC6M\Q0TaYV4AH.F
f?R8+&_^0]]aH^fINgd]AB.c6LJST&DE(1Wa@1dXW.N@&R].gNg1VP@]O&@4_9FP
cJ?9f#CX:&2@P7@<)4577B&P=_9eN[TUZEU?++CG\ICPHYB41c,;6)=@:=,.RD:V
C-05E]U\_C)AC36U4.0]],=T.VQg#LZIX6/#\V.(?M0-&PDV0R9,K\bX[/A?2a\L
<=cg_V^[(L]M59=gbBI_=1^:&U@9\Dd7(,H?(4ZU/7()1:cJ2YI,J7>(M3b5^5gf
=R,Q;V#?MT_6O56#S7HR8PV<I;d8cdK1GWa19TC3)A@K]5@VWLM3=DWOFXZ4O:;C
8FPfL8Z_J/C<&^.B6NUb-=bdR/EX.XMX6+fB;7H@60/+O3)2()gN?aKc\9Lb6F[U
B^c;SJ&QNdL@S(7F4MJ^JRg6I2B.S._=FVdGA]NHEFJPA,Z3;UNBY3,9S6(>?Qd#
c;=8)&VcI&NJCB;ALbT@c5D^H5&>1R5c/3ES/N:S?A_LM.dM6M?S@bRK(Y=7#D(N
5#.U3XYNfO[E?&]9=a>O)N\,OVeLQH;S55S,#&+X(<R7#7@3<U\SSb,9gJX2.3>]
N;;&g-;>PR)]KC.eM>6EXF7.Y(e=_c#5ITHIeL&X<)OIF3XF90-PEaA)f7SFKf6O
YXK4C8:[_f?T?#^2FMEUDP4@W/]DJB^59RZ_K/.LOH[V3La]Tc77-)gEV??6F@g?
c\dCJ8e1<KU)aXN:&@aAbIb&=U6f^SD/.@bF=PX>(+eV7f)>8EZe(41T3a+Ye>Y5
3_B_Z&e5_c1C\BWJBUDD;bF2X[(aCF-:bE]K/gNB4.U):>BK(U.XSSA_8Q9#O82G
GbAVO77?&._-:?@=HH<,0T(5^N[+15(>&ba-9+=PY4UH#XH?(-0+ORY@W(9.Me.>
g)H:3<1@PYL7fg5.c6S?LfB;[T[D4/cKTe1a6;[<B4#5&Uf3CGeWN3fFJX#0F0e.
CQ#(e7/Q<IBGa214HVbcg1P.R8+J(I>YQIBTAT>&HEF@=bS/UOGL3&7NR7,1;N[Y
4[Z\fANU+?XA/-J;e6U2O?G)H;bF7.VBEKf;8X+8]E_gJ,6EVce2dA4?HRZX)@.R
c:29BbIHJ(O@B;IHH_U/:_JH[V1@\,OLe8+CdN5FY;P))9C=Q<G?g_[PY+a3DN#M
L,JYAZJA63FY8T0Z_HD2EO=Zf&Q,8]+4Q<2^TE]@\&>Cb59C;GZZ:[8/VMR,V^bZ
(Oe1?K@gNMcLI6:;U>_gdL+;>(Va&HL,#T>.=K3&F8>0:OJ)L+d-dX-,F,,WP@40
Q#LXV+N-_DM4VASfGT=I@CLVON8C49,.6]Ub0YW&NQTaZ2LKZ-\d(\Z.Ga2J[LJ&
^[HJ^NM0?B^bVLT&LT[g@53SMK./#L#DAg)WB<2LE[LVEdE2BNT8BLL+:0<8g76D
TM,E&2EK/\D6)Y+B?<_4+J]1I3IQ/&];CB+4]&S]7Pd6eTP6fZ41F8\\.(0EL+b+
TS<51=]2FX2ZGO/VE>>6T5XA?[^a&Q7P?c@Gd?/7WU+=-f4D@I#YZ/:5b=5YQ_K_
6(>)(VbSM(dXX(9-bE/fQ:\4/\(C;#f;VK>#80?QBN9O9_g_B1:[M_0@#VRB:LB5
L_>]-bA\V_N6S)@SRL_?R(/46E+,ccF(N#5BLgI9D#2b^g[@V/Y#H<.]caD97(IW
2\RETccbMaSCeOHJ@T+OZ:OI/b4X#Z+=GZ,0&6a[a9?fa4]/N9LADUB2e&3HZJPJ
U5=Kf;)ATE#N=aI&(2#Q/RZ-2fX+>@JcIC@?1A,<Q4^9,VL0+fG@U2]I2ag[)b,A
?bTS\1)0/JK/E<&JMbgb2NK^NG\E323RF]6@)57CKYb78.M5XCWW(dTEH-<<T+Mc
)W:A;[&VMd.\PBD6fPPEgD?Z]<2X6[MEJ;F/I?.E/HQ2f_TcM&g-,M,>^]B[L4M.
A?)a(_X4LNQ6==S2#.;?YgJMI_;.9LKc,Pb,ITgdcWLM<W#8L;Wc.YNA7U869UZC
1MLY?ZV.g2N14?/:#5PE[[R5[HJ72:a4Pbb6#TXAUP_b(WQVA,.-&.<c6g)TJZ&&
:g<a/P,:<__4_X-c<V[?=3_/;04T2()c2fV8TO@ccE^Q/W6&T@4X..3.VQQDN3U,
BY0X;db0fSQ.7\3XOTD2EL^V(C^b.F,R>K7HdFL;#E2(6N=IeccY(+IB\63;X1dF
4.Qe(@S]=QVZE3gY3;E4295(9XDK<YCO&c;,ZO5+JRRHPdB4aaD^[+AYY=#4:PFL
V+<JZ)b_3T-[-C^)D2Wc9IaY.4_d)g&D&)Sd_^dZ>f,OZQ-M[3cO>6?FI[^G1c\R
e[FIW6PM&ZEBf[I&MFCT/FVJMbOR4@5R_0O4Cf7(/OTJg?0U/RDV9W+1YS.Z8[J_
R@:=:)?5-:UN_@S#/\06fVb8JA5HZO380Z(G0(/\8\TOOT;+8[bDNO)C@(GWS3Y0
@;:O:^>#3P4gM+.QGAT#-bX[(0Y)H_CVT_?^8.,d6[<-WDVeYNLL1@I9U5Tb5Ob#
ZK^gH<[gM)C2cV/EVa=L+fRGN1SKQS:++&?[ULFN\[H37J9Q9e<MQcfUd754/.J9
EA(e\B)W>KHLYFVD9IJMW1aFb-FJ3dM>9C8gSN=,5XF7R8-M[B-;RZ_LR#4eX(/K
?<V<[.26b;Ua#(J#eP+>MO&/P1,<eS_6L[L7f;,EX;P/<N9ZGP=Q3\@SE[G2U2-:
f.PYDP[Qe&,?>[Ad^O]^\84/,Q[GaE@O\ca#TA,GL/=/<AFEOFTXC40\,#U>,WM9
L2MO&G<JG@HD:FA8=T/(QW?XS_-#46]>[?aeF)W40G9@AIU&)(e/GA?(#BeLI/D+
FId:e4X-9#+D^9W/F:7eeK?C,c0H.(^TU+ESZ]&3X96NO=]gG2_Z8.X)Z(R]PI?S
W2J^cCE@0M>--7E7@@-LCCC-:#e@&WW#J=+;KT]/XTZ/>\HdV)^]\OMF5f=]GLgg
<><c.0@WB7[2IgA=gUc4(V]JZ19//5/WbSA40Z]8&Y(OfXRZM>4/X\<d>8[0QBX@
7><;3=;4:@D6R1c#-@f,5@GDJ#EMJN3H#-]@NcD=JQd1CCO,771.1-bL+SGf<,,L
&TV4g]KTYb8&O)UIZaYA,I\Z)Q+VLQ8J>O#DHJ4[LCS65#ZaJc0_)?G_UWC#bSUK
^-YA2;+82U\R2F/J#aCTfD0@a-6\^))JXAWP-=H8RL#07MRKSOC&SQ[9Z^+X_(g<
PO\9NdH32FMOgPO8g/&A:a<<ac45^dC7dMP;3.,91CS_?99e-SgOWbMV+R\V&F9N
f>XHTUY7M@<RDO(X-6\e:FPN.a,[ea_IY\fR@YW?5^;5W=e<KWb]<]c.b@6WSMC.
)H/Z=WJ50XT>PYJ[CB^F8FN&#DT+6a62HES&d=Y42\M=&HgV846cOX-dWZO5V,ZU
W>>8O#?+8f2H^>E+SYKD163M0a(gU-E(ObLF-7;V,);M/D86(U_\S\UWA7Q<;/)]
DC:;O.L.M52YI?gJb1AL?6XD/D@D]>aW#[c;?=c.>CQ[H_FR@D/7]IC++6G]BeA/
ST\-ed2T<FQKD7G+]8g(/^dZN1Z4KARN7dL#R.^;&TY_-5_QR)7Y9#RQ6YAB7<Y0
XYN1GQ5C2T9I1H@GP0#@(#8>;<W+,L/6E;P5&QJ?L&/L5&_dMR=Q42A]+GFO,MI7
;fD6991/<D9..-6cQU+;3DAYPPBUSZb]ZO3GQY7<R3b)LP.<+=H+>P6Fe(&_B+1f
GQD+0b+VgH#9#4=Ne)/1eW\\D;F6NOJ6Y8?S#,NG@E233dVK#,];@QJFLL#AaI>e
Y@>+T6^32\[7XJKN;/(JG4UUAZBTc,+\c7;;UZE3K.ZDA8caJXa7Y=NIU<9>6\UB
1,d0T;][#cLP/5>K\SVMd[[@^14S.5[V9G:>d\?,]G-66,)UZaN?].NX7V6(\(\H
ZZ3&SA(?LN(^J6UW;=\I^5N;IG_SMMUdBRg@(cQHfX]2BM]&&B<^TIIGFN2AJ73)
])H?@B@&.f+NUQ3?SZ6.BKTLT&R>#a.VI\3)-#6g)>]2P3P_F/30,dNb_,Y02)VA
ILEcFKgP=?&ZXPE4;E&\2>:aIQg&_(TN4?[F_2G=NS5e)(:PaYUJMK4dW44XX2E=
^>DR#G4L#b+_I67Q/FNbc3.BR:7?.&N?gPa7L6Fa&F3-EUSG7g-K4_CP^#?dSND+
UBX\4FP9?QCR\2DB#fGOQa8Le[ZW)[fI=#,,N,?Q.2QEK\39KPGBJS12>Dde.<(;
)P9-HR:^VU0a1RAc6\d(VY,VV5FAfG@[;<adE3GRP/TGGMONI/=d_:M=K0BL2T,L
<+H[G.5:HT8HB6H+TE/M;#12-4Rg?7\cEIcJC\FTDeg5d<=Nc]0cdZG7?4Rc=/.&
.IAHa5WI7Na7227;;(Bd_<BN6?M,8VRe8^91SAV.CBIG6@#&;.G;[Q)OGGR#OdWQ
213,M=(@?Lfg-CTcO9\QI4/f=N6M\7UB.&&6AB9^BDa&MaS.933gW6),R?S]Ef0X
Kf;_fZY2L#4PgfAg[f\aPH]IXOEW2VEC.)LILOU8B(^M=D&-UJ)9HE^TS1OL?VE5
S(Qe+3Ub5L\9_\b&Wd@:XOSf-)OQ2fAR9Y+U4@J9d8O?Y9g;.1LF=E[9RTc^&Ya3
/4aD-4Pe(<D-V8aaVC>-S_RCDKb6\D,ULL82)gZdB/(&SI7A)E@Z9U73F4##&,b6
KWCfG3;F>=Y9M,TA9eY3N&.8H_cA>XO5,.O/Sb?-I@I/fCFC[6AM>_.7T@EJ6g>O
?^P3a(bIWb8<Y<-3M;@,(\Agd)7JI7Q,[cV#W?V98,27)+MJ(VHX_]dLF<SLV^b9
4PJ_UE=NZXb6/8RT>cX9BH>9,@?Y0WJaIDTM[&?O&FP&1GgC(dMAQbddP0<.P(N6
5O+RO6XLJ1QIB,2@)Dc/QRBKC9cREg>KTaET-OLVF[\XQ;ABD,NfHgOJ3.Y]K03f
4a>350_^Q\(R@F=ZFKO/G>5P>0Ye2\DH\UXE-51W]V2H9cUOIYQZ+FKJ3\;8UC8+
OJTa\2.>dQ4cWd;T2[BYPfP1X>T[@/^FG)B<2819Z8UR-_BWQ5.TJ@&7:GP\VgV_
0g8&?I.,BHNdQ?ZD34;81dA)NUQA#_T53D2PY(BP>IKg2],S/cdaRGFc\XEY4]-3
aIO1/(\3T15UOAHR49fJ-WV&1Sg6>?S4b?a]5NN3CS?EBVVf&UV<O-UYNJAL29C]
Z5,]<C-TbR?4E__8Y2B-.COXT8DY8eCMa7#?@6@MP>>CaJb84Y[T.aA&;-U<9NX)
GcWWKD5-OecVV)bLf4_TM5AVBc(-DZ;&?RQ]B2I-BTX22L@_bSH)HfJR#@8BMP6Y
,,W_/S3eYWD0L3_4C&Y7J^fH0EdW,81.#4:8LY&XQ#W-#YV[_]HgHG7A6,4f@22M
7cD61[\P:@]bDVNTDe>I@S6E_S?E4BCWYA=S)2ce(&O0F)(^JTH1))?QOdeVdMd)
Z/>W]Q),\b7.6]+#.V:B69LIC\IT5,+=.Q#PN6R[S3D8_=.[,?,aMKS&ce5M4FJO
MI8e4#[f.[a[R=OVb/VP[7YfK4W-JFS30^\?GWV=1Q>G,A7,M.3^A#WIS,agMNYQ
2:,ZDa&+218W=AGda(MS8M(f2=GaZ/edd;#g\6O[JH^Q6(,9DSGA&QO?QfZJYa4d
:dN3=[6\6O7/C:DA=&5WXU,@:3#PA1YEA_F?EEHPK]+>RI<5)ZA:#3b1/S0P:QVV
UC&>21Fcg.GG+^]9_(N<3.AF/\a_==OF)-HFFNeT:8T,N_Jg<<GITJB(0b=8-33S
cI3K6=XM?^LI>T;e0=)D](_-1.b@OaK-L8TA&D>28a0M?-e+Y;QgR91?PG.)RZPV
<6-XQ7^E_AGHYNAR?>RQN/1,^0D>gQM,G@L(B=HADJ(39db&bfEJZIc96KY9_]Vb
5#G6;0=8PfBUX\?>2V41.QKe]1-CY^_4V/ea<QH<T6JV9YN+g4<,W#fLXgNfHO4F
ICD,UET<<BS\dE3-D]:?aP8&3PR_--YYIeZ8TGMROA[Z17dY;\6DS4e6>YA2L59_
8@5/(Q/dV]\KT?P1D<I8E9.A\J=K_(/E)cAD[]]D0X)FE\c(LaPB,&F23S[Ef35)
\YJ>S+Q7S2N10UHU&,a?02&@@#DU<FRU:+<@#D1OfN.>O+bZCfR+Wd(3+bO5b_IP
\MPJW4WY7eK2bM^^^dG<?]-gG7cW8;U-fXC(-5I;N20P6?)J?M#6Z@F^<T^8UM+b
SCJ30O(3\:f]U.E<^[3/_;dAXS1#_,#BaU&P;SKb71VJ#=]._/&/F+Z3FJ;g5#eW
<VNX\WP5LNdPU2N.K,^M,T_b17EW,0_64W=Ref@fG]+GWALNTGKJ]YF0C([@KE>f
)IU3f7VH]V_8<O6VIcf@8^_J1bJDHR;Z^)82Y&a?g/DCWZ\e@T\:CG4R^&.XdM).
0TW/fOc0=Z;[G.]:(#4I5K?<HNeXa.c@W;e/3]<C4dXY)E@Tb]b;aHb:6&G7(DK[
::JCc9-3)N\;gEcH#4,eN^N^Z-E=@V&PMK8:J])]BRLXK#&UE\XgNS>I-JVR1UAd
D/_5N8]S=+H<P)S.I+N)c9@2d;f+JJ>.=Z;=^@(C2gb;]QMc<cL0Y-^G&1)^,Bg>
Z#RL4VL+^Wg8Ee3=IUFa]9f]M^?a,d>WEOSNK#NfU_)C0PL-R_57IK.KO>_5H_VT
?C1FLJYJ\2D8RXc?7NI45B_T27LRUH\UGK-<Q=IG30=(T1:6(5CeI;_?\c4W.d=a
.OL:O8Yf3)NY(N-:F1\?0=Q3WT?8&bV:eO,N,aZ7BW5eCLB<aERILY04):;TB(NS
Ra;J01WM,Q,MB#9K](QgHN>P\1=f>=1dE:cb6AeLVI3cOQ+VV]^:Re1WC2JBST_+
>\XZ&c#:?U;3F)YU.W=R6+<)?RbD\)\-CGIN\SP(_V4)XNHFSSa6NDC6fI,L4OeP
.NUWSZBS2/19@R7\eS1a4GF^S^H].SJOWbO]@670[G=6UZJPGCefOPMNDF=:]9IG
bS:;YSQ9G&W_Bg0TQ2AE(UdY@]-A3R;INZ3[13_5+R6.SPT2]5X7[?Ee>AVdRYA3
M/fbZ1A_Z_d3VT2_6Z;gFH+8fO=+>_g4C^OXG)+@\5J00c>fcYQSQ_dQ7X>7bI\)
4>DdRQZ.6Z?8C[;eIDe,f#X7^\OZX41UC^,-b@D06?D>1NB5[Saf<\>6-NRfG?2a
eT\GaFR\I>BQ=QQ-aMcf+,F1B@6@fQ)9F[?R;Y1?+R@Af/[X/<6RQ#E4@DV+LeLG
FT^/M#M?aL;2SSS-G87#@BFZIAcdg.aFDaJ7OgLV1-^0egW\)P[Y9R;UeR0gXGSN
YaF5UORGCCc:@::LOd69#<T]-^-&_BAV4,U<3BZ,/CDYcdA]4V3dQ91BcbRa.)KN
dC.U:Q6b+;QJ=U_2DX\4\7\>Od[eGYV5JY&NIdJ=R>NEJ@EV#XeVUM@?9@0ef#4[
0?[5^3.R2ZLAVC;IDTfRQ9GEDY.g7HH3ZD.,7gRX-2WL6UZ1HKO?DXHgD0[/@Y#T
_aN[Bg.\28.1Q?;D4I+fWA@#P<WbX<2I9A7\Q<Hg5OAIg4A^O79P,N]e&E@3(<S)
KC1(+BB]eB^QR9++gL7G)KYQ7D0+7^,?Y;AXI5UGZ&Z@N#^K0U/5@@)TX?Nd37XX
>A/B3g>^7M20<MQ017E-J<L=IQA./4:;#PQ_#MEJQf(VL&?RB]S@Ib055:\:D8a?
LBF3Ea^9.A_8^BI,PLed>IE#K8CM/,>f8R0DV-/JL4c^HC=)4S&HHOH,KR+H5\VI
\;^LYI^(I@Y.7T>@a&O.SN&</PU=?>-./W,dU4^U/X]f/=R?5_6W=-B@WO+CS/@E
9Q#8MX-,HbaNfJgBe7+?G53/;2=S>JC_J]:><X+EH@EWHFe;.VaJ#I+^=XB-cdBG
a_F=f>Rd(.HS5LODV-)QK#P@P7/[G7WO9._,A(Re.=6);T1#(>F>F2&^ceB_UM+<
@aXBe?JV2+EcOG9LC\5\Q0NT605R.:RWf1d>HG>RP&&Z53Q[K2[b:(2&A,\:Ka]2
Z5/U9L-TZBV(CR2_AM6_c,1V^fL+^P4F;b_)be&A@A(I],Y1M;AF&:/e:dX9C,#_
\PbMQX?5(Z;;+-&,X[E,QE;W8PQP_LKbdD39#>eLR4)-^4G_^?8RE.?[\XeJR<ED
DT#)?>0#/>bI#S8D[)SG^N#>Oc6DU.^0\ZHK^:&]^+I:e-I8)7ffGY2O9aPV_]S^
5<JRU5PHQ4-E\eMCfZB04ILfB@Y2,>/A07()K#S.NFPH9<&<6RGZcY8NK#E;X-,8
>SF0+2U.P47Z:^;Ia89W)2R=,A<.e1b\>?b</WZL7\]&a8DNfO>dRLVS<Z;BY-8G
6,_5)-)P:WOJ3T0[&+-HcV\fO<\2g#74.R<W4:3N#Hf#Sd.WTKEWV^.K2T^+_HP:
8KR\70:@c#g/7U)b/\F(U_+TS^(bSdg3M8=\[@NE,A3M/(,TMfIO@84T7_TQ_Q_&
J07LKU4T?0LD@G(W]RQN;Z@/9a\XBTdCU9f]bWAcMMCQR?#&96JX)1FS69FM\(>@
aQLM-.49K/[K.f@P]:#ZP)8EYeKg,UXYHQ/95H8c_UO^_&WU49_aQ@]YE-8HbWV^
0.;FE\b0(2;?/H\7D1U9H#=M,]5:\-^ZA>7f0]?bK/N(SU:ES1ag8SK_=S]aTW[5
Rc/49=\f[g@-MN;bO6]091[E_2G5</(-aPaJ.B8USZ#+b0.3QJ_@;\JgGU3AI1/&
V&^/CR0+ZF+87U<M6)Z96FQA1HfEH+(4Z=.Kab@5N3MbT.\LG/2O,g0<Y4_-Y-8Q
Gf;1526>Xg=IGfA,A+]QP)H05EZ#c]e,=e8Fb..g&aB?-XG=J3+/1<;1,W:TQdKO
?Ta9P.]6-03573c2JaXf]S1#>5Q6gLCR;5^83MU2D2@_S6ae2eQ,D2U?TeJ1VHc4
;B]=WC-P26JEb/>O@#16b#&.QF;1UHQdZU:I-S(_8J/+@^/X61R2)M0@@Z\@9&cc
NdT_fSgD=c:PB_#3(UI</YNfaYbfe_.=-O;@\2[NF7[#S=?Fe9O,-KE=OMSJ.D^R
BF)I8&e)Y;D-cTO1,J97PF(FDXgW?7M=a01T(J\eH&LgG5(T>FRKf<UJ(E&L,2DG
WV6:FO>/B_cOUgNDc<N[5QKD-.PT;QKOKCA:)5b2FL6U:AcLaW-KHCE5:IBFG(PH
LgI/>.Z\IDLB5aT3BPMM(<K1H2(ATB3)V4W,#SPC6A_a30_T1dA7&Y]Fe4^+G<3W
c,dX?@SAHQT)/M-L#3VKHG;S&]^bB[A-CA[@(#d/86BOYdgQ;7TdG.OAYM#UET>\
88B\:N^e17]Sdf&b2Uf_2f@>eEV5If,\:?O9&>gI?J^d=]e6?FI8=]W+H?ENO<E\
=.M#b9/1ZFDV<O]-+=7K(/W:^^:C7;32+@IcT],4/]?ga1N&NcS:AN1#b@DVc<,M
GTUE]QY:ZU:.R]Gc6RZTJUaNY;Tg:d;G,<]AYXR>]bOLG>A4bNMYJC_:#[QOZ.X=
P&L3F4(17+F/:FH>UHaS9H8H7\_dYKFJ+VFDZVBGN6U7_<\GBZH(fH,e]2W@?;@b
NY@MO0--JRNQXI#U)4YG5.O8;=We@W]]#eVB#(cZcD_3Z;8\[g-C@60K7\e[(-Qa
=)_e]SX#eA4CPOJa??N2^A]+d/Q6SL^4-,\f\b)))b.d@H:;R<TS:HaU(Tb,NJHX
C61^.K>/#:9f>U1205H\L#:6+&g6^>bE7#S2-dQZH6aI3TZIUMF7LWRN#_@&L_H.
Eb&KD<adB]cA\XGI.MaeFXYT:NH#:BS:O.Q4(&=F3H=5]&/+>>#^)f-DKKN=)1\&
f(/P7;+1WQ4RTSGe5:bL>1PR#MM8(+eH3:-gAQTL\;c-S71#Lf:dHJe_XeCEbbI3
(7d1I:UF1^I8G4#J<59#SHVGaE@4GVAB#,1b\DN@JPbGSR4X;P#3f.L;gKNL-EZF
Q@1PYDKRe\=TG(,5JRdM-BI=DDCS==Q8JY,Bd_Bd&/3VH=Jb.(06YVYc_a>c-?]B
3GQ9CP5HXPc.LIS#JN7^-<9:@]O:@6-&S1^^DJ:[-GR.GQ<<dV^8V0#N[2J[K:9Z
LFT<&F7RUUB]#6KTQ:B;B0EXH#84#._KgK2FEL3]1Hg6J@4Eg4(gg\#2a<S^0W(9
R6>.SJ;\6=[(5:\W4GfB7\2#3HIH,P[T,1e-KL_2>JT+V;(E-.4@f0KXfIJ:SeR5
C8BKQ6Z_ORQbVOgR=+IO.@&IKDd5-U89SKdOV=f4fEc4DULKf+N2bLVA3@,#(&a/
\#Y;V^VJNE+P(K.2F_6[<AA3c:[F<?:^H6KB^E4LHGSXL@SeccKf0&P6X^BfdRG;
_UGIO/64,&Rdc<?23b/J(a#;^2(Y9PaTEVV#=b=UW1fef;\AR[3g^VH6NAddWdN)
G>2<1S82VW,YZB9WWaY:X5fa(@gO1,YBNU_#bPBd_:7.[,7HG,L8)F0](TGa)LG?
+MSI_Wc>:d)1S;_GD[LUa7<LCR5+;DZ?6cI;]gDN3==2f<7GY[b#]]^.?gUA8&eA
N6)c5RTbMC[K,O(.V<5X:f#QeX,f9=#@Ba?2H<@+fd\XLZ4a(\P#ZX4U\&RQf\N(
F&H:<\\QRNZGEFCFG/]7b,+GO1F4f2M53U;X9C:[(a@DXGSB1D/.=,GFf:\IB;,Y
c>cHDTGcX>/RG_J5Z>NN3&A\5B91KUHAG;K]M98\S)KaKUWH7K04=Ggd,I(2VaS<
gB[fd:2gaSTJ#72FN(QBAZ1V[PD1[Z/,TK[8/@R:W+-M4\UO4>#IVOKg7H14=80f
XBOfB5Q>+1835LAK/;^^93Md0&CG=S?8+?Gd)5D]=fIMKTbY;N)DaGV7RPRO,&cH
ULaK89:HL-5PX9eM>M>[Wgd2P,aVR4RYD^@6SdFM][#IFdNWa_2e^<_:GP9\f/R5
#EXJ#DC;^fH#W/Ad,+\L,@>[#9\.^TTg<\48cf/4KGYPK&+WL>^:H;:ZF?ZRRb53
P5aNEZ^,ER<A8YNZTgQ>^WZ2U=3KTC)?g<8R4(XQf,<<QN9]aYH=EQ2e&?):I8/E
04g@JQ>(P#3KD68?#c2Fa21G2AAR&_V70VQ2S5:R]F2[[>2&Z48.EaJ[6L928VSF
H;.R#==,g@?6VI<0YK<[PGUPUH93QFVa+cV\^[^H7S(01D:e@,D3F72ce=CgF+@?
^:<;aG1TLUKg3JSBFGG<c+gbWO>_)TO<B,)0F/2_8_K#E;\3.bB\</(PJ2f8AE_P
[a\#[>J-VXGT:1S:J9FG=U8&>J1218AWMO_?Qc[AV-a9VJ0SE@DY5F=&U+AJKU4F
[QLcGG_]=g8PJG35<0.\N6e8b2c\TKgQ::Yd^bQ4>)c>)-#B.C,&>B5EV((2#0fS
4U9ZY@KHD<4;ZacAR\CeZfY3-I)Cgf5+RSZP<1[[ee]CT95S0>]/Vg8=BLSYKN/B
U5<4-IO6;@XE1-0Q-C\S\0,(.+MX+ON#gX,AKAMgXSJ5_(L8&D9DXPX.S?\M@AEE
AF1[gF_(A+H7C7^J52I6ZJ<@^..))R05-#LGXNE354W8X8c4af6dG:bHR,SDE\II
f\aE#W2e^\Z4MKYXGC)1,-E9>e(:_I<V.3b43\Y9\@e&GX0Xg^6<6/+)01)_b:F9
0O+#LQKAd4)TY2Pd[K[O#DHWVR-@&]5T#Xfg(XfX2_D\9/gMFTH\D-e5e6U3.QGS
E/@6QdY5SSEE)/[Te)8;_F7KKgKecbY#1UW1_J-8ZbLBQ)ecgQ=Le_WBdd9IZOSW
@O-+G[I@Y]/U-D1>UEd</6>c-8de^4.1;(T\0_RaO@SAY-/;-8]R:KBQQ8BF+>//
)b9H?^N]e3:K]EIXI:U,J2FN:1\/cU[1<PHPgORHHX2Y:U0f\3VO;ZgD.]139CII
L..]:L6JBKL&G,=.L&<M4D65d/ag4(0(;V207(,9b<1W#Z2QQBG<(=g>CMgGD>b>
RD+a6LE)UB\O]N@<8S,V=78#.S?,0BIU1#:8WZ)XfVKU;P+Q1&eO+I;3UE)2S0,E
(;);^UJU3#Be=T6Id8WE@R:R1:1#[UZJ.>YZ;Zf-_cL7)#ERB22],[YPBAPVe65c
Ed?/91?#L-a2RAG6\b(CgB/S)5A:PF3;ZX@HZb0VWOKFSER]:KF7:)@8F<#U5W>^
+/S_GRM:U\bO_Y2(EYM?bKOP#0\DGf=+/P#7L0V1XD<,5bE>2].OP?M[+g3Q3N/S
3NW#EdL[(VV,_Gc/J,/#:8Q1:.:;P><RD?4F/J:W0e?O>Af:):Z4)DN;BbObe:&B
acF]8F8Z\5&P=5<2<(9.EeSM]b(1HOS=@</_8J:_WKOJYa1a8g;4E7&CZB3+d4K,
2R>1(HV]#g9=\75:1=\N](I?A>28.DT3,VbQ\MA;FXZ<G4?b\aS0261?)6J#P5I>
a6D1;L\cQM><HD0B@C<WJ>-R[IT:QAMCg4WX\H780FT9Ea;>S@cSDRK/<JHPe4#Q
Z<KW7<=T>AQDI(E:A-8),0X/e+0[,e2XdJ-P<XX(?87P_#b[+)]0R^]2Z:J74P0f
]660IMC4IS-M,KeYE\\T.3IS-_I1b.5(S]ZD2,I.Oc1JT3BBGC_IGg:_\f2PbEVZ
,XXa0I5[BO7=fcR1PP?8CQY?3RNTV31RK@aCeW;JA0(NO?9C;@B6-BPT7.bNSDb0
H7Da@.[]He-/I4B]:eIJGf=?@0(d83KAPK#\KRM>]9L>UdD@#P._I9c:/)L)D0fK
DeJd<M7GY48a1B-5d_A-g<ZSXeX2UUHEg3;.O?cO;b\<Z99-@)G:7+Vg;DcVL)\G
4a;<]KG+WR]4>DC(RMPdDFI_dONB6VgF0JUdF[68RPAITO0]P0>65R;(:JND=6(3
Db9H?#5;1Af<5>PZ,AI(M]37XJ,b0?4_+b_CaE2R/SP+OWXD#4dN_,+V?N#Xaa,Z
GC3SH77U@37DGd@YY=FJ-cA09>8#-bb0c^(>\+,X\YS.3c5MAHH,5F:.5QUJTCI4
Pb.2&W=Of(JIeT5JcNABT,H(ZZaAMWd,AW=?,V:QRgCR:X\M0b1C;aH>17#EYY>M
MKO,).dBV+6N=0G940,7W.V8-ZEC02RBIgf/MSDO)F0-65+#R\&3L@0eSG#cR[H@
9G1GD_SRL\T&]/I914O895@=@T/>@Qc[b(5XS4P+c0:2UN7LD/_aU;IB^3_L)MA/
8eB73+&((bL,]+@D/TS-KX+a@Q#Eg]6b&8,=b0B;eb@@_b<Ic_J-VSCU)1G#Rfc,
/E9^IW_5G+O3R1M\6T]R8MJRA=JU;7f<(E\1,G9HVFbSHZ-Y7.[eX83+PfY&PR:X
NPL<Z@c>&/Z#(;1fNf:5;9\Jd8<Xaf4QT:R;.)R\9H,#J6\:U3?+2,B(<KG<46K1
c(G(g,SfJe]SQXY_O@.+S@CN4JHU7#I2AXNRL9TS?<dC4L>U1)RgOZbLg61/F<+U
FeM/+68g&G6B;(2X_R3_X\8UKADF;a@g;a9(cSZUO#MGSUMQL(fMHBW<K335f9N#
(REJ;4[@>2ZM2;4;Y9EH^9D7UC#P9g:HL:HRCMF;g)MX6f@/eF,DXM@LQZ4U7Y(;
W6^J_]5@C6/+1Q?)8JaYD>1-G]Ef-g>01QXZa5ZG19\10;ZKM?E,>f9+<F,PY(TG
@0#D7LCZWES8RcW9Q.gMgK+(NG7+WL._-VN>Yf=^#W-1S:T&:&0F61<fH?.V@HG.
0#@&\cS6CW6DC+2c_JDT)Q2FCcU\>^@S@C]]ESW,O\(0+Q@V?Y7YeUaRWQc-K9eD
3NAU-M-BQLKY/^0=[D9I-SSVAL5c]7W_J@+dAbeUURf9IZ(V5;7R3bL?dIW=M)[7
6>bW@?J;_/?NRZOY+#AfI#IESC>.2-:3I;X&<-;8=:V,=5;d_dS6:/?&#<6;V3<A
g]E6,8A5/J1?[ANH02#5-3H2##KGA##.T[\CX[74S;I;U^Wb=dW=JT1;_4Q?e=Y+
0__b1]/U[78cVTL):<+^agZD-HF3@aaI:7(D^?(gaKbM?^O?g22UQ@J3BAac9T)T
YcIfd1fgTO(SPZ@NWDS_&-AH^B@,WY3Q+?N&#GVf/b.+\#4Gg1K#g<UcTE\IF?]X
-Q3&[;-:E?JYgdZEPcNf;)0<X[L7HC@V94(Wb=5GeK.@&V+W7VJa((<W8YWJU,J7
96DRFI;c(\>,F142L8_2RaKXHF_c2=H-Q&XH818@?[1<OYUOL.#+(7_1(B>)e^TR
5WRG?.FH[dfV29M+2E=0\G),Q@;SPO\37]C&U,U?c)E,S<d^b_C[/-G]F5U[DTO7
>>-:P4XEULJAA0D=D3(VGZN,R@X@;F.Y?#,?gcJc8b.:KTCHGbZbZB&f,dI]/VZC
>7TE:98bQHZ>^?3d[3TaST^=+.ARQ?0SFD>D;;;9IWRg(WU,c(/8PcFOAISbI22F
fP_=3ZfNN3a8F>0e[-IX5fY:6AB=KMc\OO4\(PR/(WJI+g6W]N(]IB8\eUF&19CP
X.866,9VUBa<A8@ZMcg#b9^4Q1&KLA\C7WUQD0^0C.EM_aKaK:V?S:\55#RU+5MO
<XX:bXAE+\\+RXSNJQ,7\4]d<ffTNE^B<G^X3.^:27+#=P]7_1Y0#?->C<C#;EJ,
EUcVP2(L,MF\]1Lf]67g;UT[6P-1N^49Y6EUGd19:KR]7.c<4<_?RQaaR/JB6=>6
M/8:K89EM8cWYF1:N&SP@+N/0#0-O0/J_:,dDDb(>X4ca8EV=:V57,98Z9T4O48R
Tf-Ab[#VQbK&bbFXO_Wf@TeOQ/HLE1a]&f2UJBe^VY-,.)OR0a(3&L@XdSCTUaT_
_>c+X=d?3>)@F5VX[N]DRQa??Mg2F\1O/FZcTN0TI<9I:?;UV/gVd0=V:7@/M;N4
WgR[CFI/P:B=@>gM,E(X,D1OOG@9c=bOU-4C_I^4cI2,@N64]&7aO5E34dRB]J<;
[#+&HO1][[a<TNCf^>D]aHTeE<R8<);=NRaCd-^\;V[_:[(Wb?f+\:e/f87<a->]
8Ue++>,[QF1Cb>XBB[Gd6Y_29MD\bY8A0=+#:TS:KX(=I:6IY[H#SA35]P,.&@-G
QX^OL^7K7Y^W]bZ2E827e6)V^3^#c8Md[>c1,b4Z)<E]NfS<G3X7Q/QQH7K^-,CN
Sc(.Jf=?4&f.=JeGTITg#2#W^:,N7aWU-4D/_6/?FHECHDV@9V]Z?=eRMAPfBcXc
Q/#?7[=#e0S=Q5JUR)fGM>>J;4=TACEMI3EfCGE.eWe5\K3@BPVLLD&^>K5EE?ZR
LadX7c\9_T7A2D)XCb1=FE3I8M(#LRF_X(N+E=E\,:PbF@TAV<15,fUB^I@(;g04
a_=)D:U@1g1TSUf/(]F7b)#H:gE?9dJ0.COO2E(R6cN9>ZGOG;MR\)KA9JV.0Gg.
XR])+Y7N/>eR5(OJ-?2LS]5O=SKCKN7@b/dT[V8\F47M2<Z]P\@CS3\G<e(Aa62b
_5;:?_.DBE@@J,BDU_WNf?PBW3CL)HQ<9@?&L_=&ICLKc.)a/>Qa?>9\A&<8MIa^
Q?95.d25FKX1::;EPe)VLSV+OR_/G+fBPC.X>YE;610]HE4M[69A(E.>4P)E;Raa
&a2Ka9JGDe50(=GO-IAJ[.B,I9XC^1M8H3<)TZH__>fXH50HS4)D4eQDZ/R+\.f7
)?&L81EgZUC^I72C?KH,bR,#MN>\NASfL)[;IW1KWA6=[#[_Z-Oc]?d+a39N=14E
g&0>45CNX5:YZO?FR&[P[T\XDIS^U-F4e(/K]==I-X-^X:0L9-<ES7D,,#G2I?LJ
;:&&/cJ5TW33&==L3\19]a]<-6>7:RT#Y_JHSWA-F7A41QZATPL<)_E_CcEEIdBL
POaY8\LT3L&CVX>-=(;:,A<-BQN/52NG/g@?8#;>MHD>d<@R+G0\dbC&S,007#Ld
61f_5bN(fL4e19LBBRV_9A)U7SJ@G=X[W;aab6AC4.#F=PVPV\)SH7QE-f^9FJd8
+[QU&E&\3DSgX<IVJDI#WY+-+,1)deaE,ba]>>OgW]8I3_fU:_XUR@S6RZZN0:Qe
MN<F^bC[-&T;H)-7-UFS1ZD4AORFHG_Qf4SbdICYf=K&.LP_],_D2H>J)LKS#d<U
MWBg8(7f5@T8.D.<>YG\f@Sc1CK_BO??+dDd9MaXG(gXBXC34X[N>D3TL@P=>K)+
,WQ.\GTH^MgGH9Mf)d5eTCP\KCM,0=[.=;]DVXFc4(HI6Q[W8>XGHJ5#0H5&,bOS
SI@CQM4G1WKUA7d;<:0fe3@E&M49>cSYH;6FV0/Z9Y<3Yad4?0V-[WGd,-\EL#MN
>#I8^.SQ2:@7YgbG4ff7.2K,ZIXeRbY[I_Y+,YU-a6>]0][P/3OPX<>0C+=>cG9;
MGBG94F9-4TR2A,DJSXOIQT]\8^,Lg_6R20dLZA?DDSJDCXKD>HfL/,cMAG4:(,9
a;JC:0#CG,WaCT:dI3d_<[.+fBJCL:/CJS)=,;b[5[#D73G2<Y6=V=EB.cadL,Id
S1GP+&BIUdGJ+^9g(+g+3\4gZW-P4:^G[23SaTWX#3.05CSgbLF#M>f3g,#^BMJO
B\6MC:EQcQ\?Y-F</\M^GC#ccC_O6eC/W^5.B+=;N\>\/?T\<>7-^3Z.VD[=X9O1
?Nb6G^-344eEbZ978^fLC;U/+_<G[.CNFGK6<^SR+b(3EQ+c;+Z^GNST0GTNC^[(
X2g?P/G&UNRgJUdJHN2Y6V=XS7IE?3)Rc2G=U>&c)?\J[cTA)/YUeX]M+YAWae\O
GW4/dJ4CG1=1(/\-/?PQeKAC&I)>[=-E5JAXAN?DM+.gCHCZcE?]>CB>&;IM#]22
X60DD6[?_6[K@_,VL#BNa]B<A14a5?VVA6?1b[[(WNTUK,ae<_GMDM\;-c+XO-?-
73-51VZ5RD>1?MWS:-d)K0/FKY0[F>YB#NDW?+@@F0BM>40&60;].ag<GC8(8AI/
C6_4V[K]Zf3.eeM.8?KYCR5&IV3Q,U8EZ5b(JPB)K>gZME=K&_7.YC5XU83D3,Tf
QVKV/Wb(V[+,.FUN3MU9gBQM6KfaaN_a1.?^4gbDR0NZ,,1cRa3PgZH(K^\T3TcW
K<-K\.3LK5W8Hb&/_GP.FA/MNCS]H>H9=<30J1.N6THI0B+gPN8Pf^[<:B5WTLY?
9/6Zd@5ad-T.\WcH<OJ,Sg&797#fRZ82&JVPDFFX?IUN&H>+#SI.1g71(XcZ]S4X
QAABWXeLA4gOg3?UPb4;\C>a@]Q\6;4:c,TX5C6X3H54\0;#:cJ<XWI3fJE;QI+X
(MP6]<^c?dcgQD/Y.KRWf\f7;/;G/50WW/&=30&<(XJ7OcG&Ke2UBVYM(9@fJU07
Z,fb\3cC=AJ6Taf\]Y+9I^H#KT,T\2f=BBIUK-ZR[9fcV.(?F1-E.66KK]R+?AV.
PNUb<C2g@RLV9E(-RVL>^VCEL<5QaN0/&d10T]+A]H>TN[.#WgV<DHK/7O11W>M-
V;;a29eH#P<;C]U10B.GDaA#129DR9c2L7X@I]K[9B2D;X732V0[]g@_;M2NcVgH
J>#5@-D4&^c5TgKE.+:(CV4g)50^e-CfS;YXH3A@X]AOGO6SBSNQH&0.KN,@.6^J
=3>\1G<KD0P>.2<J@XU7_b_Lf,+b/+/0ffc-ObC=(c>gWbef0,3b@+MQ_4QWa4A@
0RDV7f]W&WfdCYe5P1DG9Y;.4gc8gJ[Z<a8-1H5<_QT/eJ@8ABa.QXReFD(T=@Gd
AI)03^J/?BcAMf,,aaFX_YT+#P,.J9?U5EFW(YPgL>cW7:EVT2M/C6>?6#-.524+
g0C2]5bAfWZ<FDV(,Z:\JKKXaWJc08:RD1?[:2M\[HI_J#/;N<HVS]O&a9M[I2?/
N<e[5)_19;X>[4,\5AX<cJM7JeU++3W376B^,MESZ@eHbSgBE7f+X_3O8WG62>9V
73=U67/,\(63f_BC[0C)+-4g1C^#2[/PZIT-TbAb-X9T?_eY2_X_>@EBg/-B(NFc
FQ6D/+LbH0aM81E1KS?bDVeJ,1PF7;]>ZS7TB;#/TLN1YX&.-aI_K\.6FQ,H,Y0U
STX2Y@08O@cCTPKRV2&75)2EC,A2N9[0g7Z[]=aAH^]W0f?.e3OX)d3ZMW?7K1-R
Ef;ZA1GVbK+;92MZcg\ZY8EXP];VMaWUa8UNS>X[W9<_:OW#B>>8DT&e<\#M2FBT
/Ha<LEMSO/aTUI+\O<,@g[cO4Gb&3YbO9^5CQ>Q,]J_&cQ;>WYW(X6Y<79=C(GS7
WGIGG(=9C.c;6]+FaHa?cTW6K>bg)?RC8e6/^Ge/#UK/97e@V&OSc4]QI3IfJSMO
.WfXJGJ3:7K^S]NMM\+,:KCD+ETg2SW/I\E=a5)cI@2e&.2A>_[VFe\PM?#TN>Xd
Kd=88OceCK92G\.J42?U[0LPPR(@Sbf=2M4/:Z)D5<\C4<cMb&A8=+E(14#T?262
34MSGWJX5\UZ_(\9PF19##<Sg7O.C;6I0eAFTL4E/aSP)AS.?f9BN,N=eF14:H^8
5F=6bAS:Z:?/[V8\eW;B_YDd;A&WRX[62=@G-c)98\Ic@_2J?dZ1E\dffDbQZVDB
O>e#\@.F84D>?eUg.GP((GDX_@M2)8&?d&1&\<7<HFPe.g58^C:,2[VHDBH&#(LC
D]J<V5S2H4<WQEDJZA>AMN+#f,NOUS#4H(W8B)dQ;[,g=0aQ[bSG#PEY<-8P4V4,
g.#NKQBZXU1@4WdJ=cA0^_<Ybg8DLPB#P/^PNVGS-BMYC35\Z)OQ5R;7A@3P/S5>
+3Y.CSUTfN.84LL_CK?[G[c7AZWUPfP+>aF?0\4.?^.ZcV</GQ+0e_9A&f9+/0)S
eF7JV(BQIS9[R)Wb11B?eQ8RROe3@B0B@SI+RO[K+()aQM2H?--P@#4Ia?IW(68b
XR?[[Aa;]U@>TFO#-(L.[e>VLc_dRWS\_:L8>7e4/dQ^>]<22ZdBNd9.&&8>AF6<
2Peg<R\eD2\HOTaC5c^b9#,^b5<=D+&C9O(T)W:Mf51,YH6QD80IH[1A^5Z&f-@P
W&\b<OZaI/)IV=2FT)X76(@T+#34<JU/9W[)@TWL,T=?=+a<<e8,3ZL0LA8[NF:M
2K40;676YR;GD6]I(ZQS+B3bYILd#R(ITR=:V1H:,.EF#W84--5O^K57B7)@4-S<
7YDfK7/L-04WHd4W>J+^@TTO1[[RPJN)7V[J(c]JdD\OQ4\:M]dW(RD4=C7M77)f
WgG[I);a=/XJDRDc?L@,e7I@ePWLI54I6bT+-SK@g,R>ONHf-D9@a1_ML6L<63)a
I?7P0E:.L#AFJ/CfZ7H[aX+W3A2YNKcgDM9R#2HLFJ@J,?O^+3?AX<7ZbJ59TXF9
42e(&+RGKD_Ff6+)9LAdJUTJS#a&5C2GIa]G1GL_cY(U/KTC1g\;(QOA/GZO#d4#
^/50Y7Y:0ObWJNfP?IVfWB6YT<fdA\Q[4-+8RA@@,:aOG)PgO,G.QZgEOUce\Q1D
GSVOF@a^ED77\Ue+3[PdEZ:^cZY6e0<I:.H3O^I^[MHac6cD)g4;\-\9[TRC\57Q
]CR#_&>Y/8YR#bb:@_[NVQBG,@UcSG,1(IeGU[+e[2O+cD0R=B8a_KAP4<:I/DG4
])I?V&g7GRebK:?#I(&/Le?7g=F)1WdD(\5I9\:,7Zf3@QND@;4V/S]e0&Y3EA3b
L#@D03/H2+K#JSZ<LET6\Yg43GM0bW8T:73@8]<:(6.J+)3AdYW,H;&<CJ89N&C\
J&^3TCN0^OAQ7KTTG5(^9(=YKBfd)aUVK176c)Z/=Z1[VFQCJ[(bdQ<SgI#aW1_5
HDeU-7f+b/185bD5I;KU3(V5,5Egb/QZ@Vg)D&,Vb]ENL]Mg5,]QU4SB<0e]?)D0
.==UA)_J(IV@M=LPUFWK+1D?^.N@>+S49ZMTK#R7/N#)8K979gU(SJZ8XSE]0a](
6a4g-?fG3Kg5D,Hc6AV6NU0QdY]41_=g28GP^-&HUbNa#R(^0EG_JN@LX31N6JQ9
9E#+c0IR]HNe@F#<ECACD26>>O&MKHU0.c\#Q4IROENJGD.bF9[0E?EJ>1W=6N/U
&9_ZA\+.(d?E,@/MW.IWb(M6Q&UGA(Tc/d/C4][ED+NgK2R<R,ebP3PWO7H@4>;W
0I&+5g@UYOUgMfKb8F3.P[)f(d6HX:GG=NTFM,Zb[SC)c1MYDK;[KI:bM>^5O,K>
FF44AdK#>[MNZMM)VBM=2/#Z/=fR0\GWYdI^W3990_WVbJ(,?cH63>T)#9NO,5Je
TW&:4D&aBC/K=V.1)_-T-5b_ZC,.fA4Y74)^,-:[Q;03/dBW9N+JFA0AT@UOVWg<
<#N[=,4?RTIcI0;T7BgGeHO;6)]C6?KOJH45]BT,W0893>OY\JeZY?I7(>57J\f<
1?K2<1+C-/V[JM:IMH,5b)V2Q[E16fG&P2Rf?Vd,cfP,K(L=>A-Y:JFL6O51QRYE
K47&/+<_bZ).J@dB/(?9[VP;7RHT.>H16=)\IU@9ZgRfcW+3X-_7Sf:#f[9/8dfQ
J&Q1O-Sd\ZdKV6Ocf=8H>,7:#3SG>R^bNdMQ.ZJAJU;a#F<&_g2Qaf;UH):M.2LH
W-R0)F6C+9H5fc2XQB5OGAI=.RK4Pf(9_9NO,9#=F74OX2U2._590RU1e?2&e;RZ
7gGBX_5R/?A7N<GU]2g?1U-(H-6P]&N5dQ/MYD)((=-WP(e-H0be\C6J0/;NbEc?
A#5PF>..>bU?11G7SL+<fDc]T9Z>1Y9PY]:_+Q;(<ga;<8f4,c>6BaaJCN#:JA;A
4S0d)3();]+e_b2PUY-Ia<N=6&9WXE0NeQV@07G,+e;+6W\J\#e>WO<Gc0]I+fA]
.N?dEG)D]:A[Y00g0X>7)Q,B+7J.;<3ca7ENU8<VE=-:2AU.T-^)&If._7#1JX>?
c[=?K&^@BFU/9LZTWJN70H<V=bQ\3QI>C.3J7:98@G1I-U(1@G2@eacS=:8>>=7H
-3C:^HfKL(L+S;+P7C<#Qd,-XHR8J09:f<_0NUG2]?-dQI[6O&L?bHT#LR;QIHTQ
.bIJ5^VGGEK@?GR^4V,G)9G6TE8Afg\X[H?WT=+aYcT=_gOX:eQ5e1RP-d/ANI4/
?dI[,NfAOL-b57(c&03OgWY;A50bC2O6F/e]0P/b8D91VW.B,]T<dH8CfDF-8_6:
ad09SE.2Z+gf\V,Z3+(&b4BZZK,=.^RZMDf(d4E3?\;3QS(2L&-Y\>N4@WQ7A\V&
Y#2^8VB2O]B-AM&F\]M1f18B96POTG5a0F=2PH4XB>Z0Z@G#O4)a3(/Q(d858IBK
X]A;H0O)1OY=F]d<(/5RLLF:;I^1<TVU/E5H6Wa+F;6CMbLOTAf6J;I,D+B67Q9F
KWZ6^_Qc9WG1a9Z9&@Z@JP(;U;Y@6\OVZE&C0Nc4#.af@A7NT:/R]>c:5G(4>V9^
Q4ZVS:JXJE08;5(6)Y,9U+94,8W9JF\8):dYXXJ#N-;d2b;Ue9cM.Nbd7/+^&Cf4
3AFA1Y7^Y@T1gWfUVRD=8.9PDLdf#<5-YcETN(<Xa8=5^]gHYX84C4(b[]9<BVM7
#PP]2A.TX3H&(3Q8S7:=E>QOf(ML>AUIV9UY@(-G3,.&f9K4cIVdQDN0@4XQ]JbM
_R:8C+@7N/7PM3N)54_;W/J_@[VebGDZSL8QRT^:Og38JV,D8UII.TAP_a5bDN-6
2E?J-Y6c1@XF1;_2dB=H@KKT3-[;f7R9XOdM>@<OGL31/@T(#F^?JL]FIO0BP/-7
]=O5\G_N0DORB27bGT/+(N=J1e5c[AS01=]cX.(0ZaZDQ+E3GRH?XX6>Q#1,Z#=b
0DE(f+@/X9,YTg4VN&D-d\Y;,J\C]gGU)WA6:O]W(FIJ_6bLFGDI##ITd5H9F6>S
XB=+7?g[eXLNS#YS/8Jd.N3@)P1JdP6W;HN=dLR8;_]/DB.:HAdHF^UaA;[][L9A
<;XY;Q].,(fJ>)PaGfS69ATGceb;ScC29H@ZIfVVDR_Mf->5f+^fFTBMXI[1/8=g
Z&(EMF<>=I[MUbCBd;Ff[BB/M]f8\?C3KYO8)_<2/O:V7#[)A\d2XVd4A>a^CL@)
0;+D)TXcV.KL2X(_,1\gPTA=bXT2+dSN5BUNZfL_B<CX0+DFJG^2BBFG^[E6K><R
5\-LJP^QcS\[FF#X-6_@D4O,b/XDeRKdIVWX=4\1]B)EL:]aCc>F26L_EJgZa,:f
KMb33@^OcNd/JL?^UV&Rg^UNB<U1U=[]Z4)f<M8A-7MMD]8W6>0?ECIGA6@(OP#g
&AEJ,d\c:<[dEXD3/7ROD84+Iga]GXUM4aG5?8QCfS;T.XfF[7LW)X4)4eF(IXJT
7>ZNS-9dVM0feY#>:[,=7Nd0PH_@B/AFCHIK_0d_R;(8Xf9K4=bY.P73-JK=GE9_
X#_TO6?Y#f=Te[c39a6)aGfOeKJ/VQXa_<:LOVO?e29;(/DX]DOW[?H/9)DY^5CO
DR1+(GFU2K5_\@LR,abQeP;IF>V7O0PH[?VJNO13U9eaGBD9)g=FOF3eYPbgB<ec
P;?<Zf1,]3@2,f_3+91[M==5##2^XUZ]b^;\cDa@#&M<X;^^+AY=P+e].PQXJHZA
5Y#L19SXM^GfFT&_(TR[ILK#b&R?TKN6;M/HTQG:H8d3UVY+M1IFEY#OeB76X5];
7C7,Q/.XRC&,<@21[e3G>G&&8EJ8Zf;\Q:fWKD#A4Z\)2U2P/UNC0R)@e;5^0C,&
X6F;+&f769A4d,EdUX]UTG,=3e;a>&\+H)9Q3+I1APD86S;cG#_;aJ;P2+PM^#:D
X(W6;<aBL;61D\G)aTg?]BTf+E2g/,6GTfgJ[X+QE,0g(X1ZZ,:B[1&O9^=f]U0,
/a?7d^O(KC>;1(e/)e--ZOJUQeKKYe,PGQ?+&J8(6O&d(P2=H6?U4Ac_f:/V(e:8
T7=(-#4feL_3PJ0OCV#FMdCS57TWZ7T7V2R2eGWcgO,VWFMA<P+(e-cRGD25T.cX
XPT@RAMfZJ>665[7?[-&5BRRJ9+;.=e[2c2XZ1&7ZJ#0f01IKOW9aaGKcN,C\D3-
JHMXBE68a7K=\K)b(#=<ZP3X>f^V^<19@#N4Y?Kc8+R]X;Y1-@c^YY8-9V+,3ET:
X-N\I2-eYA4C;]@G\2GbgH/ObE<HF,ZQ0)7g1(6:&Q/=_)0R=C:Z0Z^==),=9(=,
Hg_(O<8L?0M_/VWBbe2=+)]CBDeMGH]BH@<I2g-);)NFLNBC5BBABA5\HE;W8I\]
5:&6\7&]e7&<A[?4gC#BM;#fYDg=S^C,4?5FEYXQeQY[-X&?Q4a@g\AS/(f)8QLC
5S)W[G@7.O1)UGXV3.ec(+L;C]2HIaS/_&(I3+dO8#K>:fG&<aA1@P.Q1Q/c>/_?
Kc?Q95-Y(,<1B-?U_(P0^:G/K^fLE0fXTPDd.B_\7e<-/?9BOS#J-\(GM\)&g);Y
ZI9Q=_/FOOB@,=)gc9IE[4cg_<9O\68Vd:;[>76;P/#e_XK3?2c@(X/D+FO(->F3
WS]4E2Nb7O:44ZcJJAX[b+D]4/>](8d:bW#/<1PK5,#2Z8#JN_=25O3W-:,Z=2bZ
6E0O,Z3J<8de)c9YIAL8A5+]79MV8.H8VfcIXZQXYJgR.W^[f]=_R]I5?#2>:T::
BOf;RK:.9N2)HF#Q_Z1T\/0cCXWB9&9X:H18H/c=G7072H:<Q0e-GY;.=J@(NNC\
C#)g_J)II8.d>,4@:Uf[6Ta:>];.2U0&0O[7d\12:H@15W9/1Bd@LP17a8g7I_EP
U>a@M=d8Y)7fb1g0_e-P.3FSD\\;3J:2],8E]4Y<>?6c+V;D,?0,H^4WEZT/cD3/
VQE[Q]>?09T4./c98@@3^?]NL1+@;[LaV?YL;#94@8;SMC]9Vdb(CeDP+VBO_\\&
BdW\P@BfQ2\KF7(;],]9Z1THQ<E85:6>C]U+</J5a928-Ue3NCA07Sfg]b;L>05O
MPPVK@LB(7WLHYC_XD[eXXW)b,?WaGaH1]JW4\&PCHY.OA;&^P5+GV[JS<@Yb2f1
=3X-=1gQ]A(C0.19XRgUP<OJB\:7^FRYSYaPVdU]U:54U/+K=Ma[<A@+1;2@HR+F
\05d)^H@]P<;.#J#\YCW).J4e9GJ_W_bB:-ZGSF^:FTO,8444S==G/6:(TeLKeKg
MU8NEf=a?7QB89La-NB6XM=#]S5)Y+[a4[,9D#c/QIg]+_[a,QAcB)6GHN;U+2ET
_UOa]=U(J.(5BR_V+dW7L(cZQ(4HK3K3<TTFe=9(HW16P7^0VgJ0\>S_:47K<0)?
_]IJQ+S1F0YD8YA)TH)HdU]V,,JG#VLU72_GEbdGD/+_N2J)d<J0](]E75P,HMfc
-HIe;/=L/]^B\5L.BC,;ORa95SaL_KaF3a.;FF6JV6>Rf0CX;F/UO^WO5I_SLc,,
,?-24\d?0KCD0FcWHW[J3.;,O5?.GVT,R0\-ITPC2&Y^L2F-fLW>DOTCT:E[\U&<
dAD6IG?@>(3U@9#WV)#_QG)OGIJ=[0-dfH]OC\W^1V#c>5aN#V46,;GSN6Ia(/)S
M>VGX-XC0,T72CRY1Qg4<LOJfIDP]Mc//\.OeJ>MS(HR92N?D53gH4(VR\FFd>(5
6V.>1.T^+(Z?aNWI@T4>]O]5KW5.(RC:?e48TLN0.gG#0K5Sf4G?@@T93\R[1TbF
80]LA2LHAW?<T@87=5@80JX&;_)@XZ/=LVT:\Q5-RbfVD_,D]:YPPN:efEADP29d
FT-3fVZUM]8)F=O^:g>:(N@6X5+6e[f#ND0M)g7g4S]3.QP<MdJMMG&QU,PMW-Na
J4PdFFe:M9BfSK7U)P4BG4-R\5cL1J?-PNLNYUF?KK+J=ag:T?(WdJ:Z;1:9a3,H
#JP@b+A(L4)/5GT#\(_0\,3._+[,,27VV_N,E9[XJ+FR+4X236:(FBBFAS.@^@B=
KJ8beF:,c+M13\N@#_4g+V+O)9H6#b:V^U+_Z[QQ+IYVE&8+a.9RYV<4KT;47QPP
@,^AH]R?b-^PB^H-(#:d&?d=?/7L_YQX7S>GI40,@A@;R[YVJ,X6K9,]RcG2:303
V3M8(DDB^F<6I:DSFK4GT>A:\,CHRJ[2\dT>J9H=+14F2P1B8><82^JdR5((5e&S
9_>7>F[2HUf>KOI[bHRZb8_ERT:#O=N+@38U0T6M_V;,Y-.Oa;0feO?4S&e/4;\_
]5IC3I4R@,JMVc/&8=4;4UP=EbcVS,YWS4c^GC[X[G]JNYC#[?[5S9TYDSM;ZMe/
ce>B]/I?7]<+6Y/8+FR[5f^]P;95A3<A6DZ6\G1(SFMO;JZ+XIQ3HK,T_.?@[^.\
PQ4AX6BU6\[\9J5T[JB,)c0D&S9.^BCI=423VED<baU,_S]ef55202UGTJ\LB5LF
2<_ZODg(771c@S>8]]d6\]RSU+=AHf(^4f[^.5Z]Jc9FPRXQf03g#g?&IA2d@@:4
UCBW4K^2\V<Q+BF30Hg91KZU)W3]aFfYeSH#L3670\ZCc_@0>Df6#1[Qg4/U6aJ4
@,+=c:9+&b+ZTe5<c38^J[W.8eaGd@DCD3B1[7>J50^/CMU]+8agS1[]Q6V#1SV&
^M7R>3E3;A=O4<2#Md;B9e.T.65H=FE&PUH<^-IH(8WJBT2EGR=&_PD,P&VI?JI:
BEF-eXR\g3A&KDS=K]MT\ZRCBb/\-H-\;W2-KQGXBNgQ[+^LPPPXI#6?XKE^Q5Sd
WZMU]7[78TZ,<XbbI^8YVU#Od.H(29T&#HLE,814f/^C90gVCG<IgC8-W?Y-K,4_
UQR@:I;ZaDa]YYQ^,#4T<;[A:eb1M=EP9GET7O(<FD(]IW.&U0bIP>]/IGGab=Ra
cba3UA[NL<1Z557/6f1\66UN0VQ8&>HJR.Hd&MeY0ZQD4f\T1RW/@XI&P\?_GgC4
ggeZF20EPLO2ZO)E@&Za,cdJ-+QScb+[T_>CY(70W4U2BEY@SB_,[^,-D@Q9S@b<
&M\JaFI:;RdIgPEO#Aa3]dQB+=U;BDVdB;67=[.GcgO9ebc84VD4bOE^]4N\Qb?P
:cO[10VA(TXNZ,GF5g]8ISBH3T[)7O/<=#+Y\[?\37@+#Z41dNBf:agX2<WGB)-d
NgP(XQ-(d4cP7f9=,FaYG\cb)+GW>b+HMeWL>74G]]W)6>=OIdDM#O7XMQAC<O5c
0\Q,N7JXFB)7a5aE28&<c(EO.<@_69;,?&RY.8;W7e]CNY=eHVX=:L1-Gc>c)R)a
SeKCCH?,\/(5I3,+7;-#g=#-Z8B,DR<([?QG58\:IULVQCUS<M60>Eg\5RCITY4#
M/H5@2:D@cP=+Y=d@.<EJAGC9,f_(0D7Q8dKGS]YN&b[db4.BSN&I1H8\UI3MZL^
OA\Z9_Tc,XFQ[R@W]&T5A.N\Wa21KaaNBIENQA9e(Z);d\G/KQWUeW2RI[7Z;I/d
N[6(0]Y?D.=dN/0R+,B9VE,YXCYEN\B1UN?8aQMY:^6AX?U0)CeUJ3W(DH5D\NI2
=^c2+g-dWa/OD&7L\LbLFMLe0_EV.55g5_/QWMVafMJPAd3&08WNJ9ZW<RTNOe+,
,1_2H>H.f,U,4CEPJMD9&KXI/8/b&\.<f/3(7_#)eA1fZ3RM>#>)E;B@9H&04#:C
Sf80Te&&)B?E:YS&6C:de8;XgHZF5a+\KR/9^95gM+[4f,7aXPX7Td<Pd-4@gC?H
@]&I>ZbDaKK-C1XXZ=QEg:.@e^HI2b<,Za\I@E=U_8CZ\2eK_ER>&a?&D26]U](L
_8<P.dBDeCX<=?-=8F-Z2JGLCQR6:BRAH)T8GVW(OTE7>eXV=8YYg=TJS?YT0UQ=
&RGg4R9>;@c1&6PD<@:FMCg=1MCTbPX(L0U.NgRSYNFU2Z-JZF3<LaBg:;X;51(-
:aP_FXR:36D)R?f7CcK2g.6OU&:6(0J:@E2,LG=^=;P38.O:(PJ1ZRKO13#[^fLb
ZF?<e=bGOFJ#LSB?9CDPXdZXaCIP.B5IOM896ge^X<GMV:)<c5GO9Q.^2BJ1g>H9
7]OW<]Z5FV(761NJ@:ZH^YHC_1T_QU1Pc4U[&(W#Ob_-H0?0)77B@2;geId4a\CK
C,bcI13E&94595>>TRSc#.)e_-FWe(6.]:Y8]\^J)_]9VZE+39U=\@JF0\;ccNFX
80Q=f0;V_0;g]\^CD6D?+N<e#;[cF)7DC?_3AZQ/5DUBEJ#RN5H>VG<Y2(+T++3g
^SP7^DG<dePI]B,J@W?7;.b10+>AG65AVJM]Z4V04SR0cfK<20^5:_?4cc;fCZgY
bA=4/YV]d&<M9UYRV&:A_E#GTR.XK<eZ+b:&[]Y)&QG#UUE][C5N,OLR=K]LS<^#
;FN)4J.8W)/8+<R291b/^\C47#B5&#8cL27Z@b8@\)Q<U1W8VS7f(eN=a[.,^7e2
<=f@6=V-9Sa;W4)XMQ]\/Wb<)/<D)S^B82.X2F#eB;1M@6]HG:(HC,PFY6Z09DN6
[6MCQ,YP)=ZN6R81>/8,QTHaB^bbXMXe-]F[C-DNNKgR1dac.FS)1g=,L77f#K[9
;T[VRX<N&,9TH#3:<5/M:->/BX8=E5c:QgfI\7F57CQN)/OD4(d)-A&&[N&L-0bG
81_86IYXK8F<2_ZR1cHP\31[fZC8(\ec;:H05:.76\_YbVe3:-QH_:LTX@&D9J.4
,L_4,[CEN0LV^PNHLSf.Q[>;),@7D1Sc=OC]C<Y.]_U2I992LPU5-WD</VEHI)eg
CbSXJ/H3A9&MO+J.^(eWeDG#dOP0fSHK8>Y8B7B]TIMOMe/1?HCP),S;M_7K:?Pc
;89TdXG3-b#e8Q>;N>2/,ZA4N47ZDNH0?KC&PZe(3K7IKQ\NbF=VGKUM^JTH5I,B
>L2[,Q&fg5348T6I^-fV8f.D,H-^J@+a\0VZY;+6Xe7I2WH@2T=7.^)F:Of/C]=;
0,P,#,bE>d--Oab7@Y[>DO&>4\<F3X,WHUO@&IMDTZfG[1@2F<,8RU:GcQT6G2<,
-aUF]KA@CG[0=<R94eBb58?,]&[8?,[LAdCZ&,[9]#4>(9YTWB<4J).?2+O3;2;b
&VV/ceCd4V:F4Y2KSZba&PY.3R[25<TCbAC(=5,MNf:Gb)M&4ZFT[#^Af@g?>gMe
6^YFCH[Pf8eFd/LZ^IP9Ge^)SY_ReC>,10E[&5MU.:=f7C/(]gXNCKf1WUH(&\<8
8WM=N0ffHGC(Ucb0__=5,8=3KaJ2d:?8J5U9>61@Hd.3fPU\N7-[=OZ9fK&9MK;?
CD<5I2F<M[)ZH77U]]aX=77c?d&2b3@?+@,IV;LP1#GPGa3HE:\7E5DEDgGBa7-(
,&bBC<bYdd@V(V/KB>8S1e<g=U64JVVD^N,(M54Xa/d)@V,GD:UXfS&N6ePW,)CZ
&f;a;U4Q)]>N=g>ON679@dD(PQfHd;0g>Vc/C^]8e#/-P31f@69@&;S=((fF6gJ,
D26W66<E,=DI6bFQcM#-Qd54MPG(H&3O//GPSZ5?RBL+01V@84Z7T)GB6;CR[DBb
SJ4Yg4I30^Q/<Z.L=W76XU6b?2;R7-9eP=TTQ6gg>,<6E/.=7IO#/V1ZZ@>]Kc5M
E;A3R)c3[ZCQ9I=gbPM<)9UQb8@5AaO][S[VKDSeU0DEP;+F9G:;9-g7M41VW\OF
LH2>1a=bK6;Mf-^HeI8^9_:P.<7PI2;0&Hd.>:cScE6ED@=+IAT/;OBFLIRBSVTe
9cS8QCS3[6X?3GfbRP2>Mg>]F59>2[#-g_-cUR,/,[#:INI[E)XP]gOW4PAM9IQI
TA5BJb.WdK,VZ/O]UQLUdJ[?HW5TMJf?H6gO18R#T3X2;LOMY9JYEW3H:=D-48AF
ISd_K5>cNK]c=,N7V37S3JaP5&\)A&1?c++7,?8De24V\(U/BT-d&#bCV=]<M_FU
VU/&9(OU?#3C+BA>W1XJ@2fLJUJMB3/BE2g1<XO@B@HAQ;1EaOg@3[>P.RKKg7C^
]9dV;0V\f4f&H&#7QeGE--g5F<EN0N@]Gc[JUA2BeALL6:B^R+:#FBg?)Ef^J-.&
8JTfSa8[IdPJJ?C0F88.#ROE5_\ZT@?I=$
`endprotected
endmodule
