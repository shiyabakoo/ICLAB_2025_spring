/RAID2/COURSE/2025_Spring/iclab/iclab023/Final_Project_2025/04_MEM/SUMA180_256X16.lef