/RAID2/COURSE/BackUp/2023_Spring/iclab/iclabta01/Lab10_TA_file_25S/TA_PATTERN.sv