# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : MID_SRAM.v
#       Words            : 128
#       Bits             : 128
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2025/04/13 13:50:35
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO MID_SRAM.v
CLASS BLOCK ;
FOREIGN MID_SRAM.v 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 1899.060 BY 176.400 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 1897.940 164.980 1899.060 168.220 ;
  LAYER ME3 ;
  RECT 1897.940 164.980 1899.060 168.220 ;
  LAYER ME2 ;
  RECT 1897.940 164.980 1899.060 168.220 ;
  LAYER ME1 ;
  RECT 1897.940 164.980 1899.060 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 125.780 1899.060 129.020 ;
  LAYER ME3 ;
  RECT 1897.940 125.780 1899.060 129.020 ;
  LAYER ME2 ;
  RECT 1897.940 125.780 1899.060 129.020 ;
  LAYER ME1 ;
  RECT 1897.940 125.780 1899.060 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 117.940 1899.060 121.180 ;
  LAYER ME3 ;
  RECT 1897.940 117.940 1899.060 121.180 ;
  LAYER ME2 ;
  RECT 1897.940 117.940 1899.060 121.180 ;
  LAYER ME1 ;
  RECT 1897.940 117.940 1899.060 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 110.100 1899.060 113.340 ;
  LAYER ME3 ;
  RECT 1897.940 110.100 1899.060 113.340 ;
  LAYER ME2 ;
  RECT 1897.940 110.100 1899.060 113.340 ;
  LAYER ME1 ;
  RECT 1897.940 110.100 1899.060 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 102.260 1899.060 105.500 ;
  LAYER ME3 ;
  RECT 1897.940 102.260 1899.060 105.500 ;
  LAYER ME2 ;
  RECT 1897.940 102.260 1899.060 105.500 ;
  LAYER ME1 ;
  RECT 1897.940 102.260 1899.060 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 94.420 1899.060 97.660 ;
  LAYER ME3 ;
  RECT 1897.940 94.420 1899.060 97.660 ;
  LAYER ME2 ;
  RECT 1897.940 94.420 1899.060 97.660 ;
  LAYER ME1 ;
  RECT 1897.940 94.420 1899.060 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 86.580 1899.060 89.820 ;
  LAYER ME3 ;
  RECT 1897.940 86.580 1899.060 89.820 ;
  LAYER ME2 ;
  RECT 1897.940 86.580 1899.060 89.820 ;
  LAYER ME1 ;
  RECT 1897.940 86.580 1899.060 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 47.380 1899.060 50.620 ;
  LAYER ME3 ;
  RECT 1897.940 47.380 1899.060 50.620 ;
  LAYER ME2 ;
  RECT 1897.940 47.380 1899.060 50.620 ;
  LAYER ME1 ;
  RECT 1897.940 47.380 1899.060 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 39.540 1899.060 42.780 ;
  LAYER ME3 ;
  RECT 1897.940 39.540 1899.060 42.780 ;
  LAYER ME2 ;
  RECT 1897.940 39.540 1899.060 42.780 ;
  LAYER ME1 ;
  RECT 1897.940 39.540 1899.060 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 31.700 1899.060 34.940 ;
  LAYER ME3 ;
  RECT 1897.940 31.700 1899.060 34.940 ;
  LAYER ME2 ;
  RECT 1897.940 31.700 1899.060 34.940 ;
  LAYER ME1 ;
  RECT 1897.940 31.700 1899.060 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 23.860 1899.060 27.100 ;
  LAYER ME3 ;
  RECT 1897.940 23.860 1899.060 27.100 ;
  LAYER ME2 ;
  RECT 1897.940 23.860 1899.060 27.100 ;
  LAYER ME1 ;
  RECT 1897.940 23.860 1899.060 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 16.020 1899.060 19.260 ;
  LAYER ME3 ;
  RECT 1897.940 16.020 1899.060 19.260 ;
  LAYER ME2 ;
  RECT 1897.940 16.020 1899.060 19.260 ;
  LAYER ME1 ;
  RECT 1897.940 16.020 1899.060 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 8.180 1899.060 11.420 ;
  LAYER ME3 ;
  RECT 1897.940 8.180 1899.060 11.420 ;
  LAYER ME2 ;
  RECT 1897.940 8.180 1899.060 11.420 ;
  LAYER ME1 ;
  RECT 1897.940 8.180 1899.060 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1874.040 175.280 1877.580 176.400 ;
  LAYER ME3 ;
  RECT 1874.040 175.280 1877.580 176.400 ;
  LAYER ME2 ;
  RECT 1874.040 175.280 1877.580 176.400 ;
  LAYER ME1 ;
  RECT 1874.040 175.280 1877.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1865.360 175.280 1868.900 176.400 ;
  LAYER ME3 ;
  RECT 1865.360 175.280 1868.900 176.400 ;
  LAYER ME2 ;
  RECT 1865.360 175.280 1868.900 176.400 ;
  LAYER ME1 ;
  RECT 1865.360 175.280 1868.900 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1856.680 175.280 1860.220 176.400 ;
  LAYER ME3 ;
  RECT 1856.680 175.280 1860.220 176.400 ;
  LAYER ME2 ;
  RECT 1856.680 175.280 1860.220 176.400 ;
  LAYER ME1 ;
  RECT 1856.680 175.280 1860.220 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1848.000 175.280 1851.540 176.400 ;
  LAYER ME3 ;
  RECT 1848.000 175.280 1851.540 176.400 ;
  LAYER ME2 ;
  RECT 1848.000 175.280 1851.540 176.400 ;
  LAYER ME1 ;
  RECT 1848.000 175.280 1851.540 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1839.320 175.280 1842.860 176.400 ;
  LAYER ME3 ;
  RECT 1839.320 175.280 1842.860 176.400 ;
  LAYER ME2 ;
  RECT 1839.320 175.280 1842.860 176.400 ;
  LAYER ME1 ;
  RECT 1839.320 175.280 1842.860 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1830.640 175.280 1834.180 176.400 ;
  LAYER ME3 ;
  RECT 1830.640 175.280 1834.180 176.400 ;
  LAYER ME2 ;
  RECT 1830.640 175.280 1834.180 176.400 ;
  LAYER ME1 ;
  RECT 1830.640 175.280 1834.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1787.240 175.280 1790.780 176.400 ;
  LAYER ME3 ;
  RECT 1787.240 175.280 1790.780 176.400 ;
  LAYER ME2 ;
  RECT 1787.240 175.280 1790.780 176.400 ;
  LAYER ME1 ;
  RECT 1787.240 175.280 1790.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1778.560 175.280 1782.100 176.400 ;
  LAYER ME3 ;
  RECT 1778.560 175.280 1782.100 176.400 ;
  LAYER ME2 ;
  RECT 1778.560 175.280 1782.100 176.400 ;
  LAYER ME1 ;
  RECT 1778.560 175.280 1782.100 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1769.880 175.280 1773.420 176.400 ;
  LAYER ME3 ;
  RECT 1769.880 175.280 1773.420 176.400 ;
  LAYER ME2 ;
  RECT 1769.880 175.280 1773.420 176.400 ;
  LAYER ME1 ;
  RECT 1769.880 175.280 1773.420 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1761.200 175.280 1764.740 176.400 ;
  LAYER ME3 ;
  RECT 1761.200 175.280 1764.740 176.400 ;
  LAYER ME2 ;
  RECT 1761.200 175.280 1764.740 176.400 ;
  LAYER ME1 ;
  RECT 1761.200 175.280 1764.740 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1752.520 175.280 1756.060 176.400 ;
  LAYER ME3 ;
  RECT 1752.520 175.280 1756.060 176.400 ;
  LAYER ME2 ;
  RECT 1752.520 175.280 1756.060 176.400 ;
  LAYER ME1 ;
  RECT 1752.520 175.280 1756.060 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1743.840 175.280 1747.380 176.400 ;
  LAYER ME3 ;
  RECT 1743.840 175.280 1747.380 176.400 ;
  LAYER ME2 ;
  RECT 1743.840 175.280 1747.380 176.400 ;
  LAYER ME1 ;
  RECT 1743.840 175.280 1747.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1700.440 175.280 1703.980 176.400 ;
  LAYER ME3 ;
  RECT 1700.440 175.280 1703.980 176.400 ;
  LAYER ME2 ;
  RECT 1700.440 175.280 1703.980 176.400 ;
  LAYER ME1 ;
  RECT 1700.440 175.280 1703.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1691.760 175.280 1695.300 176.400 ;
  LAYER ME3 ;
  RECT 1691.760 175.280 1695.300 176.400 ;
  LAYER ME2 ;
  RECT 1691.760 175.280 1695.300 176.400 ;
  LAYER ME1 ;
  RECT 1691.760 175.280 1695.300 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1683.080 175.280 1686.620 176.400 ;
  LAYER ME3 ;
  RECT 1683.080 175.280 1686.620 176.400 ;
  LAYER ME2 ;
  RECT 1683.080 175.280 1686.620 176.400 ;
  LAYER ME1 ;
  RECT 1683.080 175.280 1686.620 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1674.400 175.280 1677.940 176.400 ;
  LAYER ME3 ;
  RECT 1674.400 175.280 1677.940 176.400 ;
  LAYER ME2 ;
  RECT 1674.400 175.280 1677.940 176.400 ;
  LAYER ME1 ;
  RECT 1674.400 175.280 1677.940 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1665.720 175.280 1669.260 176.400 ;
  LAYER ME3 ;
  RECT 1665.720 175.280 1669.260 176.400 ;
  LAYER ME2 ;
  RECT 1665.720 175.280 1669.260 176.400 ;
  LAYER ME1 ;
  RECT 1665.720 175.280 1669.260 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1657.040 175.280 1660.580 176.400 ;
  LAYER ME3 ;
  RECT 1657.040 175.280 1660.580 176.400 ;
  LAYER ME2 ;
  RECT 1657.040 175.280 1660.580 176.400 ;
  LAYER ME1 ;
  RECT 1657.040 175.280 1660.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1613.640 175.280 1617.180 176.400 ;
  LAYER ME3 ;
  RECT 1613.640 175.280 1617.180 176.400 ;
  LAYER ME2 ;
  RECT 1613.640 175.280 1617.180 176.400 ;
  LAYER ME1 ;
  RECT 1613.640 175.280 1617.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1604.960 175.280 1608.500 176.400 ;
  LAYER ME3 ;
  RECT 1604.960 175.280 1608.500 176.400 ;
  LAYER ME2 ;
  RECT 1604.960 175.280 1608.500 176.400 ;
  LAYER ME1 ;
  RECT 1604.960 175.280 1608.500 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1596.280 175.280 1599.820 176.400 ;
  LAYER ME3 ;
  RECT 1596.280 175.280 1599.820 176.400 ;
  LAYER ME2 ;
  RECT 1596.280 175.280 1599.820 176.400 ;
  LAYER ME1 ;
  RECT 1596.280 175.280 1599.820 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1587.600 175.280 1591.140 176.400 ;
  LAYER ME3 ;
  RECT 1587.600 175.280 1591.140 176.400 ;
  LAYER ME2 ;
  RECT 1587.600 175.280 1591.140 176.400 ;
  LAYER ME1 ;
  RECT 1587.600 175.280 1591.140 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1578.920 175.280 1582.460 176.400 ;
  LAYER ME3 ;
  RECT 1578.920 175.280 1582.460 176.400 ;
  LAYER ME2 ;
  RECT 1578.920 175.280 1582.460 176.400 ;
  LAYER ME1 ;
  RECT 1578.920 175.280 1582.460 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1570.240 175.280 1573.780 176.400 ;
  LAYER ME3 ;
  RECT 1570.240 175.280 1573.780 176.400 ;
  LAYER ME2 ;
  RECT 1570.240 175.280 1573.780 176.400 ;
  LAYER ME1 ;
  RECT 1570.240 175.280 1573.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1526.840 175.280 1530.380 176.400 ;
  LAYER ME3 ;
  RECT 1526.840 175.280 1530.380 176.400 ;
  LAYER ME2 ;
  RECT 1526.840 175.280 1530.380 176.400 ;
  LAYER ME1 ;
  RECT 1526.840 175.280 1530.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1518.160 175.280 1521.700 176.400 ;
  LAYER ME3 ;
  RECT 1518.160 175.280 1521.700 176.400 ;
  LAYER ME2 ;
  RECT 1518.160 175.280 1521.700 176.400 ;
  LAYER ME1 ;
  RECT 1518.160 175.280 1521.700 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1509.480 175.280 1513.020 176.400 ;
  LAYER ME3 ;
  RECT 1509.480 175.280 1513.020 176.400 ;
  LAYER ME2 ;
  RECT 1509.480 175.280 1513.020 176.400 ;
  LAYER ME1 ;
  RECT 1509.480 175.280 1513.020 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1500.800 175.280 1504.340 176.400 ;
  LAYER ME3 ;
  RECT 1500.800 175.280 1504.340 176.400 ;
  LAYER ME2 ;
  RECT 1500.800 175.280 1504.340 176.400 ;
  LAYER ME1 ;
  RECT 1500.800 175.280 1504.340 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1492.120 175.280 1495.660 176.400 ;
  LAYER ME3 ;
  RECT 1492.120 175.280 1495.660 176.400 ;
  LAYER ME2 ;
  RECT 1492.120 175.280 1495.660 176.400 ;
  LAYER ME1 ;
  RECT 1492.120 175.280 1495.660 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1483.440 175.280 1486.980 176.400 ;
  LAYER ME3 ;
  RECT 1483.440 175.280 1486.980 176.400 ;
  LAYER ME2 ;
  RECT 1483.440 175.280 1486.980 176.400 ;
  LAYER ME1 ;
  RECT 1483.440 175.280 1486.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1440.040 175.280 1443.580 176.400 ;
  LAYER ME3 ;
  RECT 1440.040 175.280 1443.580 176.400 ;
  LAYER ME2 ;
  RECT 1440.040 175.280 1443.580 176.400 ;
  LAYER ME1 ;
  RECT 1440.040 175.280 1443.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1431.360 175.280 1434.900 176.400 ;
  LAYER ME3 ;
  RECT 1431.360 175.280 1434.900 176.400 ;
  LAYER ME2 ;
  RECT 1431.360 175.280 1434.900 176.400 ;
  LAYER ME1 ;
  RECT 1431.360 175.280 1434.900 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1422.680 175.280 1426.220 176.400 ;
  LAYER ME3 ;
  RECT 1422.680 175.280 1426.220 176.400 ;
  LAYER ME2 ;
  RECT 1422.680 175.280 1426.220 176.400 ;
  LAYER ME1 ;
  RECT 1422.680 175.280 1426.220 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1414.000 175.280 1417.540 176.400 ;
  LAYER ME3 ;
  RECT 1414.000 175.280 1417.540 176.400 ;
  LAYER ME2 ;
  RECT 1414.000 175.280 1417.540 176.400 ;
  LAYER ME1 ;
  RECT 1414.000 175.280 1417.540 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1405.320 175.280 1408.860 176.400 ;
  LAYER ME3 ;
  RECT 1405.320 175.280 1408.860 176.400 ;
  LAYER ME2 ;
  RECT 1405.320 175.280 1408.860 176.400 ;
  LAYER ME1 ;
  RECT 1405.320 175.280 1408.860 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1396.640 175.280 1400.180 176.400 ;
  LAYER ME3 ;
  RECT 1396.640 175.280 1400.180 176.400 ;
  LAYER ME2 ;
  RECT 1396.640 175.280 1400.180 176.400 ;
  LAYER ME1 ;
  RECT 1396.640 175.280 1400.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1353.240 175.280 1356.780 176.400 ;
  LAYER ME3 ;
  RECT 1353.240 175.280 1356.780 176.400 ;
  LAYER ME2 ;
  RECT 1353.240 175.280 1356.780 176.400 ;
  LAYER ME1 ;
  RECT 1353.240 175.280 1356.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1344.560 175.280 1348.100 176.400 ;
  LAYER ME3 ;
  RECT 1344.560 175.280 1348.100 176.400 ;
  LAYER ME2 ;
  RECT 1344.560 175.280 1348.100 176.400 ;
  LAYER ME1 ;
  RECT 1344.560 175.280 1348.100 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1335.880 175.280 1339.420 176.400 ;
  LAYER ME3 ;
  RECT 1335.880 175.280 1339.420 176.400 ;
  LAYER ME2 ;
  RECT 1335.880 175.280 1339.420 176.400 ;
  LAYER ME1 ;
  RECT 1335.880 175.280 1339.420 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1327.200 175.280 1330.740 176.400 ;
  LAYER ME3 ;
  RECT 1327.200 175.280 1330.740 176.400 ;
  LAYER ME2 ;
  RECT 1327.200 175.280 1330.740 176.400 ;
  LAYER ME1 ;
  RECT 1327.200 175.280 1330.740 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1318.520 175.280 1322.060 176.400 ;
  LAYER ME3 ;
  RECT 1318.520 175.280 1322.060 176.400 ;
  LAYER ME2 ;
  RECT 1318.520 175.280 1322.060 176.400 ;
  LAYER ME1 ;
  RECT 1318.520 175.280 1322.060 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1309.840 175.280 1313.380 176.400 ;
  LAYER ME3 ;
  RECT 1309.840 175.280 1313.380 176.400 ;
  LAYER ME2 ;
  RECT 1309.840 175.280 1313.380 176.400 ;
  LAYER ME1 ;
  RECT 1309.840 175.280 1313.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1266.440 175.280 1269.980 176.400 ;
  LAYER ME3 ;
  RECT 1266.440 175.280 1269.980 176.400 ;
  LAYER ME2 ;
  RECT 1266.440 175.280 1269.980 176.400 ;
  LAYER ME1 ;
  RECT 1266.440 175.280 1269.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1257.760 175.280 1261.300 176.400 ;
  LAYER ME3 ;
  RECT 1257.760 175.280 1261.300 176.400 ;
  LAYER ME2 ;
  RECT 1257.760 175.280 1261.300 176.400 ;
  LAYER ME1 ;
  RECT 1257.760 175.280 1261.300 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1249.080 175.280 1252.620 176.400 ;
  LAYER ME3 ;
  RECT 1249.080 175.280 1252.620 176.400 ;
  LAYER ME2 ;
  RECT 1249.080 175.280 1252.620 176.400 ;
  LAYER ME1 ;
  RECT 1249.080 175.280 1252.620 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1240.400 175.280 1243.940 176.400 ;
  LAYER ME3 ;
  RECT 1240.400 175.280 1243.940 176.400 ;
  LAYER ME2 ;
  RECT 1240.400 175.280 1243.940 176.400 ;
  LAYER ME1 ;
  RECT 1240.400 175.280 1243.940 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1231.720 175.280 1235.260 176.400 ;
  LAYER ME3 ;
  RECT 1231.720 175.280 1235.260 176.400 ;
  LAYER ME2 ;
  RECT 1231.720 175.280 1235.260 176.400 ;
  LAYER ME1 ;
  RECT 1231.720 175.280 1235.260 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1223.040 175.280 1226.580 176.400 ;
  LAYER ME3 ;
  RECT 1223.040 175.280 1226.580 176.400 ;
  LAYER ME2 ;
  RECT 1223.040 175.280 1226.580 176.400 ;
  LAYER ME1 ;
  RECT 1223.040 175.280 1226.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1179.640 175.280 1183.180 176.400 ;
  LAYER ME3 ;
  RECT 1179.640 175.280 1183.180 176.400 ;
  LAYER ME2 ;
  RECT 1179.640 175.280 1183.180 176.400 ;
  LAYER ME1 ;
  RECT 1179.640 175.280 1183.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1170.960 175.280 1174.500 176.400 ;
  LAYER ME3 ;
  RECT 1170.960 175.280 1174.500 176.400 ;
  LAYER ME2 ;
  RECT 1170.960 175.280 1174.500 176.400 ;
  LAYER ME1 ;
  RECT 1170.960 175.280 1174.500 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1162.280 175.280 1165.820 176.400 ;
  LAYER ME3 ;
  RECT 1162.280 175.280 1165.820 176.400 ;
  LAYER ME2 ;
  RECT 1162.280 175.280 1165.820 176.400 ;
  LAYER ME1 ;
  RECT 1162.280 175.280 1165.820 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1153.600 175.280 1157.140 176.400 ;
  LAYER ME3 ;
  RECT 1153.600 175.280 1157.140 176.400 ;
  LAYER ME2 ;
  RECT 1153.600 175.280 1157.140 176.400 ;
  LAYER ME1 ;
  RECT 1153.600 175.280 1157.140 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1144.920 175.280 1148.460 176.400 ;
  LAYER ME3 ;
  RECT 1144.920 175.280 1148.460 176.400 ;
  LAYER ME2 ;
  RECT 1144.920 175.280 1148.460 176.400 ;
  LAYER ME1 ;
  RECT 1144.920 175.280 1148.460 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1136.240 175.280 1139.780 176.400 ;
  LAYER ME3 ;
  RECT 1136.240 175.280 1139.780 176.400 ;
  LAYER ME2 ;
  RECT 1136.240 175.280 1139.780 176.400 ;
  LAYER ME1 ;
  RECT 1136.240 175.280 1139.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1092.840 175.280 1096.380 176.400 ;
  LAYER ME3 ;
  RECT 1092.840 175.280 1096.380 176.400 ;
  LAYER ME2 ;
  RECT 1092.840 175.280 1096.380 176.400 ;
  LAYER ME1 ;
  RECT 1092.840 175.280 1096.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1084.160 175.280 1087.700 176.400 ;
  LAYER ME3 ;
  RECT 1084.160 175.280 1087.700 176.400 ;
  LAYER ME2 ;
  RECT 1084.160 175.280 1087.700 176.400 ;
  LAYER ME1 ;
  RECT 1084.160 175.280 1087.700 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1075.480 175.280 1079.020 176.400 ;
  LAYER ME3 ;
  RECT 1075.480 175.280 1079.020 176.400 ;
  LAYER ME2 ;
  RECT 1075.480 175.280 1079.020 176.400 ;
  LAYER ME1 ;
  RECT 1075.480 175.280 1079.020 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1066.800 175.280 1070.340 176.400 ;
  LAYER ME3 ;
  RECT 1066.800 175.280 1070.340 176.400 ;
  LAYER ME2 ;
  RECT 1066.800 175.280 1070.340 176.400 ;
  LAYER ME1 ;
  RECT 1066.800 175.280 1070.340 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1058.120 175.280 1061.660 176.400 ;
  LAYER ME3 ;
  RECT 1058.120 175.280 1061.660 176.400 ;
  LAYER ME2 ;
  RECT 1058.120 175.280 1061.660 176.400 ;
  LAYER ME1 ;
  RECT 1058.120 175.280 1061.660 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1049.440 175.280 1052.980 176.400 ;
  LAYER ME3 ;
  RECT 1049.440 175.280 1052.980 176.400 ;
  LAYER ME2 ;
  RECT 1049.440 175.280 1052.980 176.400 ;
  LAYER ME1 ;
  RECT 1049.440 175.280 1052.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1006.040 175.280 1009.580 176.400 ;
  LAYER ME3 ;
  RECT 1006.040 175.280 1009.580 176.400 ;
  LAYER ME2 ;
  RECT 1006.040 175.280 1009.580 176.400 ;
  LAYER ME1 ;
  RECT 1006.040 175.280 1009.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 997.360 175.280 1000.900 176.400 ;
  LAYER ME3 ;
  RECT 997.360 175.280 1000.900 176.400 ;
  LAYER ME2 ;
  RECT 997.360 175.280 1000.900 176.400 ;
  LAYER ME1 ;
  RECT 997.360 175.280 1000.900 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 988.680 175.280 992.220 176.400 ;
  LAYER ME3 ;
  RECT 988.680 175.280 992.220 176.400 ;
  LAYER ME2 ;
  RECT 988.680 175.280 992.220 176.400 ;
  LAYER ME1 ;
  RECT 988.680 175.280 992.220 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 980.000 175.280 983.540 176.400 ;
  LAYER ME3 ;
  RECT 980.000 175.280 983.540 176.400 ;
  LAYER ME2 ;
  RECT 980.000 175.280 983.540 176.400 ;
  LAYER ME1 ;
  RECT 980.000 175.280 983.540 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 971.320 175.280 974.860 176.400 ;
  LAYER ME3 ;
  RECT 971.320 175.280 974.860 176.400 ;
  LAYER ME2 ;
  RECT 971.320 175.280 974.860 176.400 ;
  LAYER ME1 ;
  RECT 971.320 175.280 974.860 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 962.640 175.280 966.180 176.400 ;
  LAYER ME3 ;
  RECT 962.640 175.280 966.180 176.400 ;
  LAYER ME2 ;
  RECT 962.640 175.280 966.180 176.400 ;
  LAYER ME1 ;
  RECT 962.640 175.280 966.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 919.240 175.280 922.780 176.400 ;
  LAYER ME3 ;
  RECT 919.240 175.280 922.780 176.400 ;
  LAYER ME2 ;
  RECT 919.240 175.280 922.780 176.400 ;
  LAYER ME1 ;
  RECT 919.240 175.280 922.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 910.560 175.280 914.100 176.400 ;
  LAYER ME3 ;
  RECT 910.560 175.280 914.100 176.400 ;
  LAYER ME2 ;
  RECT 910.560 175.280 914.100 176.400 ;
  LAYER ME1 ;
  RECT 910.560 175.280 914.100 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 901.880 175.280 905.420 176.400 ;
  LAYER ME3 ;
  RECT 901.880 175.280 905.420 176.400 ;
  LAYER ME2 ;
  RECT 901.880 175.280 905.420 176.400 ;
  LAYER ME1 ;
  RECT 901.880 175.280 905.420 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 893.200 175.280 896.740 176.400 ;
  LAYER ME3 ;
  RECT 893.200 175.280 896.740 176.400 ;
  LAYER ME2 ;
  RECT 893.200 175.280 896.740 176.400 ;
  LAYER ME1 ;
  RECT 893.200 175.280 896.740 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 884.520 175.280 888.060 176.400 ;
  LAYER ME3 ;
  RECT 884.520 175.280 888.060 176.400 ;
  LAYER ME2 ;
  RECT 884.520 175.280 888.060 176.400 ;
  LAYER ME1 ;
  RECT 884.520 175.280 888.060 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 875.840 175.280 879.380 176.400 ;
  LAYER ME3 ;
  RECT 875.840 175.280 879.380 176.400 ;
  LAYER ME2 ;
  RECT 875.840 175.280 879.380 176.400 ;
  LAYER ME1 ;
  RECT 875.840 175.280 879.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 832.440 175.280 835.980 176.400 ;
  LAYER ME3 ;
  RECT 832.440 175.280 835.980 176.400 ;
  LAYER ME2 ;
  RECT 832.440 175.280 835.980 176.400 ;
  LAYER ME1 ;
  RECT 832.440 175.280 835.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 823.760 175.280 827.300 176.400 ;
  LAYER ME3 ;
  RECT 823.760 175.280 827.300 176.400 ;
  LAYER ME2 ;
  RECT 823.760 175.280 827.300 176.400 ;
  LAYER ME1 ;
  RECT 823.760 175.280 827.300 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 815.080 175.280 818.620 176.400 ;
  LAYER ME3 ;
  RECT 815.080 175.280 818.620 176.400 ;
  LAYER ME2 ;
  RECT 815.080 175.280 818.620 176.400 ;
  LAYER ME1 ;
  RECT 815.080 175.280 818.620 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 806.400 175.280 809.940 176.400 ;
  LAYER ME3 ;
  RECT 806.400 175.280 809.940 176.400 ;
  LAYER ME2 ;
  RECT 806.400 175.280 809.940 176.400 ;
  LAYER ME1 ;
  RECT 806.400 175.280 809.940 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 797.720 175.280 801.260 176.400 ;
  LAYER ME3 ;
  RECT 797.720 175.280 801.260 176.400 ;
  LAYER ME2 ;
  RECT 797.720 175.280 801.260 176.400 ;
  LAYER ME1 ;
  RECT 797.720 175.280 801.260 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 789.040 175.280 792.580 176.400 ;
  LAYER ME3 ;
  RECT 789.040 175.280 792.580 176.400 ;
  LAYER ME2 ;
  RECT 789.040 175.280 792.580 176.400 ;
  LAYER ME1 ;
  RECT 789.040 175.280 792.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 745.640 175.280 749.180 176.400 ;
  LAYER ME3 ;
  RECT 745.640 175.280 749.180 176.400 ;
  LAYER ME2 ;
  RECT 745.640 175.280 749.180 176.400 ;
  LAYER ME1 ;
  RECT 745.640 175.280 749.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 736.960 175.280 740.500 176.400 ;
  LAYER ME3 ;
  RECT 736.960 175.280 740.500 176.400 ;
  LAYER ME2 ;
  RECT 736.960 175.280 740.500 176.400 ;
  LAYER ME1 ;
  RECT 736.960 175.280 740.500 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 728.280 175.280 731.820 176.400 ;
  LAYER ME3 ;
  RECT 728.280 175.280 731.820 176.400 ;
  LAYER ME2 ;
  RECT 728.280 175.280 731.820 176.400 ;
  LAYER ME1 ;
  RECT 728.280 175.280 731.820 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 719.600 175.280 723.140 176.400 ;
  LAYER ME3 ;
  RECT 719.600 175.280 723.140 176.400 ;
  LAYER ME2 ;
  RECT 719.600 175.280 723.140 176.400 ;
  LAYER ME1 ;
  RECT 719.600 175.280 723.140 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 710.920 175.280 714.460 176.400 ;
  LAYER ME3 ;
  RECT 710.920 175.280 714.460 176.400 ;
  LAYER ME2 ;
  RECT 710.920 175.280 714.460 176.400 ;
  LAYER ME1 ;
  RECT 710.920 175.280 714.460 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 702.240 175.280 705.780 176.400 ;
  LAYER ME3 ;
  RECT 702.240 175.280 705.780 176.400 ;
  LAYER ME2 ;
  RECT 702.240 175.280 705.780 176.400 ;
  LAYER ME1 ;
  RECT 702.240 175.280 705.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 658.840 175.280 662.380 176.400 ;
  LAYER ME3 ;
  RECT 658.840 175.280 662.380 176.400 ;
  LAYER ME2 ;
  RECT 658.840 175.280 662.380 176.400 ;
  LAYER ME1 ;
  RECT 658.840 175.280 662.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 650.160 175.280 653.700 176.400 ;
  LAYER ME3 ;
  RECT 650.160 175.280 653.700 176.400 ;
  LAYER ME2 ;
  RECT 650.160 175.280 653.700 176.400 ;
  LAYER ME1 ;
  RECT 650.160 175.280 653.700 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 641.480 175.280 645.020 176.400 ;
  LAYER ME3 ;
  RECT 641.480 175.280 645.020 176.400 ;
  LAYER ME2 ;
  RECT 641.480 175.280 645.020 176.400 ;
  LAYER ME1 ;
  RECT 641.480 175.280 645.020 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 632.800 175.280 636.340 176.400 ;
  LAYER ME3 ;
  RECT 632.800 175.280 636.340 176.400 ;
  LAYER ME2 ;
  RECT 632.800 175.280 636.340 176.400 ;
  LAYER ME1 ;
  RECT 632.800 175.280 636.340 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 624.120 175.280 627.660 176.400 ;
  LAYER ME3 ;
  RECT 624.120 175.280 627.660 176.400 ;
  LAYER ME2 ;
  RECT 624.120 175.280 627.660 176.400 ;
  LAYER ME1 ;
  RECT 624.120 175.280 627.660 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 615.440 175.280 618.980 176.400 ;
  LAYER ME3 ;
  RECT 615.440 175.280 618.980 176.400 ;
  LAYER ME2 ;
  RECT 615.440 175.280 618.980 176.400 ;
  LAYER ME1 ;
  RECT 615.440 175.280 618.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 572.040 175.280 575.580 176.400 ;
  LAYER ME3 ;
  RECT 572.040 175.280 575.580 176.400 ;
  LAYER ME2 ;
  RECT 572.040 175.280 575.580 176.400 ;
  LAYER ME1 ;
  RECT 572.040 175.280 575.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 563.360 175.280 566.900 176.400 ;
  LAYER ME3 ;
  RECT 563.360 175.280 566.900 176.400 ;
  LAYER ME2 ;
  RECT 563.360 175.280 566.900 176.400 ;
  LAYER ME1 ;
  RECT 563.360 175.280 566.900 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 554.680 175.280 558.220 176.400 ;
  LAYER ME3 ;
  RECT 554.680 175.280 558.220 176.400 ;
  LAYER ME2 ;
  RECT 554.680 175.280 558.220 176.400 ;
  LAYER ME1 ;
  RECT 554.680 175.280 558.220 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.000 175.280 549.540 176.400 ;
  LAYER ME3 ;
  RECT 546.000 175.280 549.540 176.400 ;
  LAYER ME2 ;
  RECT 546.000 175.280 549.540 176.400 ;
  LAYER ME1 ;
  RECT 546.000 175.280 549.540 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.320 175.280 540.860 176.400 ;
  LAYER ME3 ;
  RECT 537.320 175.280 540.860 176.400 ;
  LAYER ME2 ;
  RECT 537.320 175.280 540.860 176.400 ;
  LAYER ME1 ;
  RECT 537.320 175.280 540.860 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.640 175.280 532.180 176.400 ;
  LAYER ME3 ;
  RECT 528.640 175.280 532.180 176.400 ;
  LAYER ME2 ;
  RECT 528.640 175.280 532.180 176.400 ;
  LAYER ME1 ;
  RECT 528.640 175.280 532.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.240 175.280 488.780 176.400 ;
  LAYER ME3 ;
  RECT 485.240 175.280 488.780 176.400 ;
  LAYER ME2 ;
  RECT 485.240 175.280 488.780 176.400 ;
  LAYER ME1 ;
  RECT 485.240 175.280 488.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.560 175.280 480.100 176.400 ;
  LAYER ME3 ;
  RECT 476.560 175.280 480.100 176.400 ;
  LAYER ME2 ;
  RECT 476.560 175.280 480.100 176.400 ;
  LAYER ME1 ;
  RECT 476.560 175.280 480.100 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.880 175.280 471.420 176.400 ;
  LAYER ME3 ;
  RECT 467.880 175.280 471.420 176.400 ;
  LAYER ME2 ;
  RECT 467.880 175.280 471.420 176.400 ;
  LAYER ME1 ;
  RECT 467.880 175.280 471.420 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.200 175.280 462.740 176.400 ;
  LAYER ME3 ;
  RECT 459.200 175.280 462.740 176.400 ;
  LAYER ME2 ;
  RECT 459.200 175.280 462.740 176.400 ;
  LAYER ME1 ;
  RECT 459.200 175.280 462.740 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.520 175.280 454.060 176.400 ;
  LAYER ME3 ;
  RECT 450.520 175.280 454.060 176.400 ;
  LAYER ME2 ;
  RECT 450.520 175.280 454.060 176.400 ;
  LAYER ME1 ;
  RECT 450.520 175.280 454.060 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.840 175.280 445.380 176.400 ;
  LAYER ME3 ;
  RECT 441.840 175.280 445.380 176.400 ;
  LAYER ME2 ;
  RECT 441.840 175.280 445.380 176.400 ;
  LAYER ME1 ;
  RECT 441.840 175.280 445.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.440 175.280 401.980 176.400 ;
  LAYER ME3 ;
  RECT 398.440 175.280 401.980 176.400 ;
  LAYER ME2 ;
  RECT 398.440 175.280 401.980 176.400 ;
  LAYER ME1 ;
  RECT 398.440 175.280 401.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.760 175.280 393.300 176.400 ;
  LAYER ME3 ;
  RECT 389.760 175.280 393.300 176.400 ;
  LAYER ME2 ;
  RECT 389.760 175.280 393.300 176.400 ;
  LAYER ME1 ;
  RECT 389.760 175.280 393.300 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.080 175.280 384.620 176.400 ;
  LAYER ME3 ;
  RECT 381.080 175.280 384.620 176.400 ;
  LAYER ME2 ;
  RECT 381.080 175.280 384.620 176.400 ;
  LAYER ME1 ;
  RECT 381.080 175.280 384.620 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.400 175.280 375.940 176.400 ;
  LAYER ME3 ;
  RECT 372.400 175.280 375.940 176.400 ;
  LAYER ME2 ;
  RECT 372.400 175.280 375.940 176.400 ;
  LAYER ME1 ;
  RECT 372.400 175.280 375.940 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 175.280 367.260 176.400 ;
  LAYER ME3 ;
  RECT 363.720 175.280 367.260 176.400 ;
  LAYER ME2 ;
  RECT 363.720 175.280 367.260 176.400 ;
  LAYER ME1 ;
  RECT 363.720 175.280 367.260 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.040 175.280 358.580 176.400 ;
  LAYER ME3 ;
  RECT 355.040 175.280 358.580 176.400 ;
  LAYER ME2 ;
  RECT 355.040 175.280 358.580 176.400 ;
  LAYER ME1 ;
  RECT 355.040 175.280 358.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 175.280 315.180 176.400 ;
  LAYER ME3 ;
  RECT 311.640 175.280 315.180 176.400 ;
  LAYER ME2 ;
  RECT 311.640 175.280 315.180 176.400 ;
  LAYER ME1 ;
  RECT 311.640 175.280 315.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 175.280 306.500 176.400 ;
  LAYER ME3 ;
  RECT 302.960 175.280 306.500 176.400 ;
  LAYER ME2 ;
  RECT 302.960 175.280 306.500 176.400 ;
  LAYER ME1 ;
  RECT 302.960 175.280 306.500 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 175.280 297.820 176.400 ;
  LAYER ME3 ;
  RECT 294.280 175.280 297.820 176.400 ;
  LAYER ME2 ;
  RECT 294.280 175.280 297.820 176.400 ;
  LAYER ME1 ;
  RECT 294.280 175.280 297.820 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 175.280 289.140 176.400 ;
  LAYER ME3 ;
  RECT 285.600 175.280 289.140 176.400 ;
  LAYER ME2 ;
  RECT 285.600 175.280 289.140 176.400 ;
  LAYER ME1 ;
  RECT 285.600 175.280 289.140 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 175.280 280.460 176.400 ;
  LAYER ME3 ;
  RECT 276.920 175.280 280.460 176.400 ;
  LAYER ME2 ;
  RECT 276.920 175.280 280.460 176.400 ;
  LAYER ME1 ;
  RECT 276.920 175.280 280.460 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 175.280 271.780 176.400 ;
  LAYER ME3 ;
  RECT 268.240 175.280 271.780 176.400 ;
  LAYER ME2 ;
  RECT 268.240 175.280 271.780 176.400 ;
  LAYER ME1 ;
  RECT 268.240 175.280 271.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 175.280 228.380 176.400 ;
  LAYER ME3 ;
  RECT 224.840 175.280 228.380 176.400 ;
  LAYER ME2 ;
  RECT 224.840 175.280 228.380 176.400 ;
  LAYER ME1 ;
  RECT 224.840 175.280 228.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 175.280 219.700 176.400 ;
  LAYER ME3 ;
  RECT 216.160 175.280 219.700 176.400 ;
  LAYER ME2 ;
  RECT 216.160 175.280 219.700 176.400 ;
  LAYER ME1 ;
  RECT 216.160 175.280 219.700 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 175.280 211.020 176.400 ;
  LAYER ME3 ;
  RECT 207.480 175.280 211.020 176.400 ;
  LAYER ME2 ;
  RECT 207.480 175.280 211.020 176.400 ;
  LAYER ME1 ;
  RECT 207.480 175.280 211.020 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 175.280 202.340 176.400 ;
  LAYER ME3 ;
  RECT 198.800 175.280 202.340 176.400 ;
  LAYER ME2 ;
  RECT 198.800 175.280 202.340 176.400 ;
  LAYER ME1 ;
  RECT 198.800 175.280 202.340 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 175.280 193.660 176.400 ;
  LAYER ME3 ;
  RECT 190.120 175.280 193.660 176.400 ;
  LAYER ME2 ;
  RECT 190.120 175.280 193.660 176.400 ;
  LAYER ME1 ;
  RECT 190.120 175.280 193.660 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 175.280 184.980 176.400 ;
  LAYER ME3 ;
  RECT 181.440 175.280 184.980 176.400 ;
  LAYER ME2 ;
  RECT 181.440 175.280 184.980 176.400 ;
  LAYER ME1 ;
  RECT 181.440 175.280 184.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 175.280 141.580 176.400 ;
  LAYER ME3 ;
  RECT 138.040 175.280 141.580 176.400 ;
  LAYER ME2 ;
  RECT 138.040 175.280 141.580 176.400 ;
  LAYER ME1 ;
  RECT 138.040 175.280 141.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 175.280 132.900 176.400 ;
  LAYER ME3 ;
  RECT 129.360 175.280 132.900 176.400 ;
  LAYER ME2 ;
  RECT 129.360 175.280 132.900 176.400 ;
  LAYER ME1 ;
  RECT 129.360 175.280 132.900 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 175.280 124.220 176.400 ;
  LAYER ME3 ;
  RECT 120.680 175.280 124.220 176.400 ;
  LAYER ME2 ;
  RECT 120.680 175.280 124.220 176.400 ;
  LAYER ME1 ;
  RECT 120.680 175.280 124.220 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 175.280 115.540 176.400 ;
  LAYER ME3 ;
  RECT 112.000 175.280 115.540 176.400 ;
  LAYER ME2 ;
  RECT 112.000 175.280 115.540 176.400 ;
  LAYER ME1 ;
  RECT 112.000 175.280 115.540 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 175.280 106.860 176.400 ;
  LAYER ME3 ;
  RECT 103.320 175.280 106.860 176.400 ;
  LAYER ME2 ;
  RECT 103.320 175.280 106.860 176.400 ;
  LAYER ME1 ;
  RECT 103.320 175.280 106.860 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 175.280 98.180 176.400 ;
  LAYER ME3 ;
  RECT 94.640 175.280 98.180 176.400 ;
  LAYER ME2 ;
  RECT 94.640 175.280 98.180 176.400 ;
  LAYER ME1 ;
  RECT 94.640 175.280 98.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 175.280 54.780 176.400 ;
  LAYER ME3 ;
  RECT 51.240 175.280 54.780 176.400 ;
  LAYER ME2 ;
  RECT 51.240 175.280 54.780 176.400 ;
  LAYER ME1 ;
  RECT 51.240 175.280 54.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 175.280 46.100 176.400 ;
  LAYER ME3 ;
  RECT 42.560 175.280 46.100 176.400 ;
  LAYER ME2 ;
  RECT 42.560 175.280 46.100 176.400 ;
  LAYER ME1 ;
  RECT 42.560 175.280 46.100 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 175.280 37.420 176.400 ;
  LAYER ME3 ;
  RECT 33.880 175.280 37.420 176.400 ;
  LAYER ME2 ;
  RECT 33.880 175.280 37.420 176.400 ;
  LAYER ME1 ;
  RECT 33.880 175.280 37.420 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 175.280 28.740 176.400 ;
  LAYER ME3 ;
  RECT 25.200 175.280 28.740 176.400 ;
  LAYER ME2 ;
  RECT 25.200 175.280 28.740 176.400 ;
  LAYER ME1 ;
  RECT 25.200 175.280 28.740 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 175.280 20.060 176.400 ;
  LAYER ME3 ;
  RECT 16.520 175.280 20.060 176.400 ;
  LAYER ME2 ;
  RECT 16.520 175.280 20.060 176.400 ;
  LAYER ME1 ;
  RECT 16.520 175.280 20.060 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 175.280 11.380 176.400 ;
  LAYER ME3 ;
  RECT 7.840 175.280 11.380 176.400 ;
  LAYER ME2 ;
  RECT 7.840 175.280 11.380 176.400 ;
  LAYER ME1 ;
  RECT 7.840 175.280 11.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1887.680 0.000 1891.220 1.120 ;
  LAYER ME3 ;
  RECT 1887.680 0.000 1891.220 1.120 ;
  LAYER ME2 ;
  RECT 1887.680 0.000 1891.220 1.120 ;
  LAYER ME1 ;
  RECT 1887.680 0.000 1891.220 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1865.980 0.000 1869.520 1.120 ;
  LAYER ME3 ;
  RECT 1865.980 0.000 1869.520 1.120 ;
  LAYER ME2 ;
  RECT 1865.980 0.000 1869.520 1.120 ;
  LAYER ME1 ;
  RECT 1865.980 0.000 1869.520 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1849.240 0.000 1852.780 1.120 ;
  LAYER ME3 ;
  RECT 1849.240 0.000 1852.780 1.120 ;
  LAYER ME2 ;
  RECT 1849.240 0.000 1852.780 1.120 ;
  LAYER ME1 ;
  RECT 1849.240 0.000 1852.780 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1822.580 0.000 1826.120 1.120 ;
  LAYER ME3 ;
  RECT 1822.580 0.000 1826.120 1.120 ;
  LAYER ME2 ;
  RECT 1822.580 0.000 1826.120 1.120 ;
  LAYER ME1 ;
  RECT 1822.580 0.000 1826.120 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1800.880 0.000 1804.420 1.120 ;
  LAYER ME3 ;
  RECT 1800.880 0.000 1804.420 1.120 ;
  LAYER ME2 ;
  RECT 1800.880 0.000 1804.420 1.120 ;
  LAYER ME1 ;
  RECT 1800.880 0.000 1804.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1688.040 0.000 1691.580 1.120 ;
  LAYER ME3 ;
  RECT 1688.040 0.000 1691.580 1.120 ;
  LAYER ME2 ;
  RECT 1688.040 0.000 1691.580 1.120 ;
  LAYER ME1 ;
  RECT 1688.040 0.000 1691.580 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1666.340 0.000 1669.880 1.120 ;
  LAYER ME3 ;
  RECT 1666.340 0.000 1669.880 1.120 ;
  LAYER ME2 ;
  RECT 1666.340 0.000 1669.880 1.120 ;
  LAYER ME1 ;
  RECT 1666.340 0.000 1669.880 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1639.680 0.000 1643.220 1.120 ;
  LAYER ME3 ;
  RECT 1639.680 0.000 1643.220 1.120 ;
  LAYER ME2 ;
  RECT 1639.680 0.000 1643.220 1.120 ;
  LAYER ME1 ;
  RECT 1639.680 0.000 1643.220 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1622.940 0.000 1626.480 1.120 ;
  LAYER ME3 ;
  RECT 1622.940 0.000 1626.480 1.120 ;
  LAYER ME2 ;
  RECT 1622.940 0.000 1626.480 1.120 ;
  LAYER ME1 ;
  RECT 1622.940 0.000 1626.480 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1596.280 0.000 1599.820 1.120 ;
  LAYER ME3 ;
  RECT 1596.280 0.000 1599.820 1.120 ;
  LAYER ME2 ;
  RECT 1596.280 0.000 1599.820 1.120 ;
  LAYER ME1 ;
  RECT 1596.280 0.000 1599.820 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1575.200 0.000 1578.740 1.120 ;
  LAYER ME3 ;
  RECT 1575.200 0.000 1578.740 1.120 ;
  LAYER ME2 ;
  RECT 1575.200 0.000 1578.740 1.120 ;
  LAYER ME1 ;
  RECT 1575.200 0.000 1578.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1461.740 0.000 1465.280 1.120 ;
  LAYER ME3 ;
  RECT 1461.740 0.000 1465.280 1.120 ;
  LAYER ME2 ;
  RECT 1461.740 0.000 1465.280 1.120 ;
  LAYER ME1 ;
  RECT 1461.740 0.000 1465.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1440.040 0.000 1443.580 1.120 ;
  LAYER ME3 ;
  RECT 1440.040 0.000 1443.580 1.120 ;
  LAYER ME2 ;
  RECT 1440.040 0.000 1443.580 1.120 ;
  LAYER ME1 ;
  RECT 1440.040 0.000 1443.580 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1413.380 0.000 1416.920 1.120 ;
  LAYER ME3 ;
  RECT 1413.380 0.000 1416.920 1.120 ;
  LAYER ME2 ;
  RECT 1413.380 0.000 1416.920 1.120 ;
  LAYER ME1 ;
  RECT 1413.380 0.000 1416.920 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1397.260 0.000 1400.800 1.120 ;
  LAYER ME3 ;
  RECT 1397.260 0.000 1400.800 1.120 ;
  LAYER ME2 ;
  RECT 1397.260 0.000 1400.800 1.120 ;
  LAYER ME1 ;
  RECT 1397.260 0.000 1400.800 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1370.600 0.000 1374.140 1.120 ;
  LAYER ME3 ;
  RECT 1370.600 0.000 1374.140 1.120 ;
  LAYER ME2 ;
  RECT 1370.600 0.000 1374.140 1.120 ;
  LAYER ME1 ;
  RECT 1370.600 0.000 1374.140 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1348.900 0.000 1352.440 1.120 ;
  LAYER ME3 ;
  RECT 1348.900 0.000 1352.440 1.120 ;
  LAYER ME2 ;
  RECT 1348.900 0.000 1352.440 1.120 ;
  LAYER ME1 ;
  RECT 1348.900 0.000 1352.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1236.060 0.000 1239.600 1.120 ;
  LAYER ME3 ;
  RECT 1236.060 0.000 1239.600 1.120 ;
  LAYER ME2 ;
  RECT 1236.060 0.000 1239.600 1.120 ;
  LAYER ME1 ;
  RECT 1236.060 0.000 1239.600 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1214.360 0.000 1217.900 1.120 ;
  LAYER ME3 ;
  RECT 1214.360 0.000 1217.900 1.120 ;
  LAYER ME2 ;
  RECT 1214.360 0.000 1217.900 1.120 ;
  LAYER ME1 ;
  RECT 1214.360 0.000 1217.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1187.700 0.000 1191.240 1.120 ;
  LAYER ME3 ;
  RECT 1187.700 0.000 1191.240 1.120 ;
  LAYER ME2 ;
  RECT 1187.700 0.000 1191.240 1.120 ;
  LAYER ME1 ;
  RECT 1187.700 0.000 1191.240 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1170.960 0.000 1174.500 1.120 ;
  LAYER ME3 ;
  RECT 1170.960 0.000 1174.500 1.120 ;
  LAYER ME2 ;
  RECT 1170.960 0.000 1174.500 1.120 ;
  LAYER ME1 ;
  RECT 1170.960 0.000 1174.500 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1144.300 0.000 1147.840 1.120 ;
  LAYER ME3 ;
  RECT 1144.300 0.000 1147.840 1.120 ;
  LAYER ME2 ;
  RECT 1144.300 0.000 1147.840 1.120 ;
  LAYER ME1 ;
  RECT 1144.300 0.000 1147.840 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1122.600 0.000 1126.140 1.120 ;
  LAYER ME3 ;
  RECT 1122.600 0.000 1126.140 1.120 ;
  LAYER ME2 ;
  RECT 1122.600 0.000 1126.140 1.120 ;
  LAYER ME1 ;
  RECT 1122.600 0.000 1126.140 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER ME3 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER ME2 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER ME1 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 988.060 0.000 991.600 1.120 ;
  LAYER ME3 ;
  RECT 988.060 0.000 991.600 1.120 ;
  LAYER ME2 ;
  RECT 988.060 0.000 991.600 1.120 ;
  LAYER ME1 ;
  RECT 988.060 0.000 991.600 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 960.780 0.000 964.320 1.120 ;
  LAYER ME3 ;
  RECT 960.780 0.000 964.320 1.120 ;
  LAYER ME2 ;
  RECT 960.780 0.000 964.320 1.120 ;
  LAYER ME1 ;
  RECT 960.780 0.000 964.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 952.100 0.000 955.640 1.120 ;
  LAYER ME3 ;
  RECT 952.100 0.000 955.640 1.120 ;
  LAYER ME2 ;
  RECT 952.100 0.000 955.640 1.120 ;
  LAYER ME1 ;
  RECT 952.100 0.000 955.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 924.200 0.000 927.740 1.120 ;
  LAYER ME3 ;
  RECT 924.200 0.000 927.740 1.120 ;
  LAYER ME2 ;
  RECT 924.200 0.000 927.740 1.120 ;
  LAYER ME1 ;
  RECT 924.200 0.000 927.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 913.040 0.000 916.580 1.120 ;
  LAYER ME3 ;
  RECT 913.040 0.000 916.580 1.120 ;
  LAYER ME2 ;
  RECT 913.040 0.000 916.580 1.120 ;
  LAYER ME1 ;
  RECT 913.040 0.000 916.580 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 805.160 0.000 808.700 1.120 ;
  LAYER ME3 ;
  RECT 805.160 0.000 808.700 1.120 ;
  LAYER ME2 ;
  RECT 805.160 0.000 808.700 1.120 ;
  LAYER ME1 ;
  RECT 805.160 0.000 808.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 778.500 0.000 782.040 1.120 ;
  LAYER ME3 ;
  RECT 778.500 0.000 782.040 1.120 ;
  LAYER ME2 ;
  RECT 778.500 0.000 782.040 1.120 ;
  LAYER ME1 ;
  RECT 778.500 0.000 782.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER ME3 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER ME2 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER ME1 ;
  RECT 761.760 0.000 765.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER ME3 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER ME2 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER ME1 ;
  RECT 735.100 0.000 738.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER ME3 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER ME2 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER ME1 ;
  RECT 714.020 0.000 717.560 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 692.320 0.000 695.860 1.120 ;
  LAYER ME3 ;
  RECT 692.320 0.000 695.860 1.120 ;
  LAYER ME2 ;
  RECT 692.320 0.000 695.860 1.120 ;
  LAYER ME1 ;
  RECT 692.320 0.000 695.860 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER ME3 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER ME2 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER ME1 ;
  RECT 578.860 0.000 582.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER ME3 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER ME2 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER ME1 ;
  RECT 552.820 0.000 556.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME3 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME2 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME1 ;
  RECT 536.080 0.000 539.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME3 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME2 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME1 ;
  RECT 509.420 0.000 512.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER ME3 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER ME2 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER ME1 ;
  RECT 487.720 0.000 491.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME3 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME2 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME1 ;
  RECT 466.020 0.000 469.560 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME3 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME2 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME1 ;
  RECT 353.180 0.000 356.720 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER ME3 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER ME2 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER ME1 ;
  RECT 326.520 0.000 330.060 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME3 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME2 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME1 ;
  RECT 309.780 0.000 313.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 1897.940 129.700 1899.060 132.940 ;
  LAYER ME3 ;
  RECT 1897.940 129.700 1899.060 132.940 ;
  LAYER ME2 ;
  RECT 1897.940 129.700 1899.060 132.940 ;
  LAYER ME1 ;
  RECT 1897.940 129.700 1899.060 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 121.860 1899.060 125.100 ;
  LAYER ME3 ;
  RECT 1897.940 121.860 1899.060 125.100 ;
  LAYER ME2 ;
  RECT 1897.940 121.860 1899.060 125.100 ;
  LAYER ME1 ;
  RECT 1897.940 121.860 1899.060 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 114.020 1899.060 117.260 ;
  LAYER ME3 ;
  RECT 1897.940 114.020 1899.060 117.260 ;
  LAYER ME2 ;
  RECT 1897.940 114.020 1899.060 117.260 ;
  LAYER ME1 ;
  RECT 1897.940 114.020 1899.060 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 106.180 1899.060 109.420 ;
  LAYER ME3 ;
  RECT 1897.940 106.180 1899.060 109.420 ;
  LAYER ME2 ;
  RECT 1897.940 106.180 1899.060 109.420 ;
  LAYER ME1 ;
  RECT 1897.940 106.180 1899.060 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 98.340 1899.060 101.580 ;
  LAYER ME3 ;
  RECT 1897.940 98.340 1899.060 101.580 ;
  LAYER ME2 ;
  RECT 1897.940 98.340 1899.060 101.580 ;
  LAYER ME1 ;
  RECT 1897.940 98.340 1899.060 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 90.500 1899.060 93.740 ;
  LAYER ME3 ;
  RECT 1897.940 90.500 1899.060 93.740 ;
  LAYER ME2 ;
  RECT 1897.940 90.500 1899.060 93.740 ;
  LAYER ME1 ;
  RECT 1897.940 90.500 1899.060 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 51.300 1899.060 54.540 ;
  LAYER ME3 ;
  RECT 1897.940 51.300 1899.060 54.540 ;
  LAYER ME2 ;
  RECT 1897.940 51.300 1899.060 54.540 ;
  LAYER ME1 ;
  RECT 1897.940 51.300 1899.060 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 43.460 1899.060 46.700 ;
  LAYER ME3 ;
  RECT 1897.940 43.460 1899.060 46.700 ;
  LAYER ME2 ;
  RECT 1897.940 43.460 1899.060 46.700 ;
  LAYER ME1 ;
  RECT 1897.940 43.460 1899.060 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 35.620 1899.060 38.860 ;
  LAYER ME3 ;
  RECT 1897.940 35.620 1899.060 38.860 ;
  LAYER ME2 ;
  RECT 1897.940 35.620 1899.060 38.860 ;
  LAYER ME1 ;
  RECT 1897.940 35.620 1899.060 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 27.780 1899.060 31.020 ;
  LAYER ME3 ;
  RECT 1897.940 27.780 1899.060 31.020 ;
  LAYER ME2 ;
  RECT 1897.940 27.780 1899.060 31.020 ;
  LAYER ME1 ;
  RECT 1897.940 27.780 1899.060 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 19.940 1899.060 23.180 ;
  LAYER ME3 ;
  RECT 1897.940 19.940 1899.060 23.180 ;
  LAYER ME2 ;
  RECT 1897.940 19.940 1899.060 23.180 ;
  LAYER ME1 ;
  RECT 1897.940 19.940 1899.060 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1897.940 12.100 1899.060 15.340 ;
  LAYER ME3 ;
  RECT 1897.940 12.100 1899.060 15.340 ;
  LAYER ME2 ;
  RECT 1897.940 12.100 1899.060 15.340 ;
  LAYER ME1 ;
  RECT 1897.940 12.100 1899.060 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1878.380 175.280 1881.920 176.400 ;
  LAYER ME3 ;
  RECT 1878.380 175.280 1881.920 176.400 ;
  LAYER ME2 ;
  RECT 1878.380 175.280 1881.920 176.400 ;
  LAYER ME1 ;
  RECT 1878.380 175.280 1881.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1869.700 175.280 1873.240 176.400 ;
  LAYER ME3 ;
  RECT 1869.700 175.280 1873.240 176.400 ;
  LAYER ME2 ;
  RECT 1869.700 175.280 1873.240 176.400 ;
  LAYER ME1 ;
  RECT 1869.700 175.280 1873.240 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1861.020 175.280 1864.560 176.400 ;
  LAYER ME3 ;
  RECT 1861.020 175.280 1864.560 176.400 ;
  LAYER ME2 ;
  RECT 1861.020 175.280 1864.560 176.400 ;
  LAYER ME1 ;
  RECT 1861.020 175.280 1864.560 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1852.340 175.280 1855.880 176.400 ;
  LAYER ME3 ;
  RECT 1852.340 175.280 1855.880 176.400 ;
  LAYER ME2 ;
  RECT 1852.340 175.280 1855.880 176.400 ;
  LAYER ME1 ;
  RECT 1852.340 175.280 1855.880 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1843.660 175.280 1847.200 176.400 ;
  LAYER ME3 ;
  RECT 1843.660 175.280 1847.200 176.400 ;
  LAYER ME2 ;
  RECT 1843.660 175.280 1847.200 176.400 ;
  LAYER ME1 ;
  RECT 1843.660 175.280 1847.200 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1834.980 175.280 1838.520 176.400 ;
  LAYER ME3 ;
  RECT 1834.980 175.280 1838.520 176.400 ;
  LAYER ME2 ;
  RECT 1834.980 175.280 1838.520 176.400 ;
  LAYER ME1 ;
  RECT 1834.980 175.280 1838.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1791.580 175.280 1795.120 176.400 ;
  LAYER ME3 ;
  RECT 1791.580 175.280 1795.120 176.400 ;
  LAYER ME2 ;
  RECT 1791.580 175.280 1795.120 176.400 ;
  LAYER ME1 ;
  RECT 1791.580 175.280 1795.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1782.900 175.280 1786.440 176.400 ;
  LAYER ME3 ;
  RECT 1782.900 175.280 1786.440 176.400 ;
  LAYER ME2 ;
  RECT 1782.900 175.280 1786.440 176.400 ;
  LAYER ME1 ;
  RECT 1782.900 175.280 1786.440 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1774.220 175.280 1777.760 176.400 ;
  LAYER ME3 ;
  RECT 1774.220 175.280 1777.760 176.400 ;
  LAYER ME2 ;
  RECT 1774.220 175.280 1777.760 176.400 ;
  LAYER ME1 ;
  RECT 1774.220 175.280 1777.760 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1765.540 175.280 1769.080 176.400 ;
  LAYER ME3 ;
  RECT 1765.540 175.280 1769.080 176.400 ;
  LAYER ME2 ;
  RECT 1765.540 175.280 1769.080 176.400 ;
  LAYER ME1 ;
  RECT 1765.540 175.280 1769.080 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1756.860 175.280 1760.400 176.400 ;
  LAYER ME3 ;
  RECT 1756.860 175.280 1760.400 176.400 ;
  LAYER ME2 ;
  RECT 1756.860 175.280 1760.400 176.400 ;
  LAYER ME1 ;
  RECT 1756.860 175.280 1760.400 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1748.180 175.280 1751.720 176.400 ;
  LAYER ME3 ;
  RECT 1748.180 175.280 1751.720 176.400 ;
  LAYER ME2 ;
  RECT 1748.180 175.280 1751.720 176.400 ;
  LAYER ME1 ;
  RECT 1748.180 175.280 1751.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1704.780 175.280 1708.320 176.400 ;
  LAYER ME3 ;
  RECT 1704.780 175.280 1708.320 176.400 ;
  LAYER ME2 ;
  RECT 1704.780 175.280 1708.320 176.400 ;
  LAYER ME1 ;
  RECT 1704.780 175.280 1708.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1696.100 175.280 1699.640 176.400 ;
  LAYER ME3 ;
  RECT 1696.100 175.280 1699.640 176.400 ;
  LAYER ME2 ;
  RECT 1696.100 175.280 1699.640 176.400 ;
  LAYER ME1 ;
  RECT 1696.100 175.280 1699.640 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1687.420 175.280 1690.960 176.400 ;
  LAYER ME3 ;
  RECT 1687.420 175.280 1690.960 176.400 ;
  LAYER ME2 ;
  RECT 1687.420 175.280 1690.960 176.400 ;
  LAYER ME1 ;
  RECT 1687.420 175.280 1690.960 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1678.740 175.280 1682.280 176.400 ;
  LAYER ME3 ;
  RECT 1678.740 175.280 1682.280 176.400 ;
  LAYER ME2 ;
  RECT 1678.740 175.280 1682.280 176.400 ;
  LAYER ME1 ;
  RECT 1678.740 175.280 1682.280 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1670.060 175.280 1673.600 176.400 ;
  LAYER ME3 ;
  RECT 1670.060 175.280 1673.600 176.400 ;
  LAYER ME2 ;
  RECT 1670.060 175.280 1673.600 176.400 ;
  LAYER ME1 ;
  RECT 1670.060 175.280 1673.600 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1661.380 175.280 1664.920 176.400 ;
  LAYER ME3 ;
  RECT 1661.380 175.280 1664.920 176.400 ;
  LAYER ME2 ;
  RECT 1661.380 175.280 1664.920 176.400 ;
  LAYER ME1 ;
  RECT 1661.380 175.280 1664.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1617.980 175.280 1621.520 176.400 ;
  LAYER ME3 ;
  RECT 1617.980 175.280 1621.520 176.400 ;
  LAYER ME2 ;
  RECT 1617.980 175.280 1621.520 176.400 ;
  LAYER ME1 ;
  RECT 1617.980 175.280 1621.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1609.300 175.280 1612.840 176.400 ;
  LAYER ME3 ;
  RECT 1609.300 175.280 1612.840 176.400 ;
  LAYER ME2 ;
  RECT 1609.300 175.280 1612.840 176.400 ;
  LAYER ME1 ;
  RECT 1609.300 175.280 1612.840 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1600.620 175.280 1604.160 176.400 ;
  LAYER ME3 ;
  RECT 1600.620 175.280 1604.160 176.400 ;
  LAYER ME2 ;
  RECT 1600.620 175.280 1604.160 176.400 ;
  LAYER ME1 ;
  RECT 1600.620 175.280 1604.160 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1591.940 175.280 1595.480 176.400 ;
  LAYER ME3 ;
  RECT 1591.940 175.280 1595.480 176.400 ;
  LAYER ME2 ;
  RECT 1591.940 175.280 1595.480 176.400 ;
  LAYER ME1 ;
  RECT 1591.940 175.280 1595.480 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1583.260 175.280 1586.800 176.400 ;
  LAYER ME3 ;
  RECT 1583.260 175.280 1586.800 176.400 ;
  LAYER ME2 ;
  RECT 1583.260 175.280 1586.800 176.400 ;
  LAYER ME1 ;
  RECT 1583.260 175.280 1586.800 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1574.580 175.280 1578.120 176.400 ;
  LAYER ME3 ;
  RECT 1574.580 175.280 1578.120 176.400 ;
  LAYER ME2 ;
  RECT 1574.580 175.280 1578.120 176.400 ;
  LAYER ME1 ;
  RECT 1574.580 175.280 1578.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1531.180 175.280 1534.720 176.400 ;
  LAYER ME3 ;
  RECT 1531.180 175.280 1534.720 176.400 ;
  LAYER ME2 ;
  RECT 1531.180 175.280 1534.720 176.400 ;
  LAYER ME1 ;
  RECT 1531.180 175.280 1534.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1522.500 175.280 1526.040 176.400 ;
  LAYER ME3 ;
  RECT 1522.500 175.280 1526.040 176.400 ;
  LAYER ME2 ;
  RECT 1522.500 175.280 1526.040 176.400 ;
  LAYER ME1 ;
  RECT 1522.500 175.280 1526.040 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1513.820 175.280 1517.360 176.400 ;
  LAYER ME3 ;
  RECT 1513.820 175.280 1517.360 176.400 ;
  LAYER ME2 ;
  RECT 1513.820 175.280 1517.360 176.400 ;
  LAYER ME1 ;
  RECT 1513.820 175.280 1517.360 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1505.140 175.280 1508.680 176.400 ;
  LAYER ME3 ;
  RECT 1505.140 175.280 1508.680 176.400 ;
  LAYER ME2 ;
  RECT 1505.140 175.280 1508.680 176.400 ;
  LAYER ME1 ;
  RECT 1505.140 175.280 1508.680 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1496.460 175.280 1500.000 176.400 ;
  LAYER ME3 ;
  RECT 1496.460 175.280 1500.000 176.400 ;
  LAYER ME2 ;
  RECT 1496.460 175.280 1500.000 176.400 ;
  LAYER ME1 ;
  RECT 1496.460 175.280 1500.000 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1487.780 175.280 1491.320 176.400 ;
  LAYER ME3 ;
  RECT 1487.780 175.280 1491.320 176.400 ;
  LAYER ME2 ;
  RECT 1487.780 175.280 1491.320 176.400 ;
  LAYER ME1 ;
  RECT 1487.780 175.280 1491.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1444.380 175.280 1447.920 176.400 ;
  LAYER ME3 ;
  RECT 1444.380 175.280 1447.920 176.400 ;
  LAYER ME2 ;
  RECT 1444.380 175.280 1447.920 176.400 ;
  LAYER ME1 ;
  RECT 1444.380 175.280 1447.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1435.700 175.280 1439.240 176.400 ;
  LAYER ME3 ;
  RECT 1435.700 175.280 1439.240 176.400 ;
  LAYER ME2 ;
  RECT 1435.700 175.280 1439.240 176.400 ;
  LAYER ME1 ;
  RECT 1435.700 175.280 1439.240 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1427.020 175.280 1430.560 176.400 ;
  LAYER ME3 ;
  RECT 1427.020 175.280 1430.560 176.400 ;
  LAYER ME2 ;
  RECT 1427.020 175.280 1430.560 176.400 ;
  LAYER ME1 ;
  RECT 1427.020 175.280 1430.560 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1418.340 175.280 1421.880 176.400 ;
  LAYER ME3 ;
  RECT 1418.340 175.280 1421.880 176.400 ;
  LAYER ME2 ;
  RECT 1418.340 175.280 1421.880 176.400 ;
  LAYER ME1 ;
  RECT 1418.340 175.280 1421.880 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1409.660 175.280 1413.200 176.400 ;
  LAYER ME3 ;
  RECT 1409.660 175.280 1413.200 176.400 ;
  LAYER ME2 ;
  RECT 1409.660 175.280 1413.200 176.400 ;
  LAYER ME1 ;
  RECT 1409.660 175.280 1413.200 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1400.980 175.280 1404.520 176.400 ;
  LAYER ME3 ;
  RECT 1400.980 175.280 1404.520 176.400 ;
  LAYER ME2 ;
  RECT 1400.980 175.280 1404.520 176.400 ;
  LAYER ME1 ;
  RECT 1400.980 175.280 1404.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1357.580 175.280 1361.120 176.400 ;
  LAYER ME3 ;
  RECT 1357.580 175.280 1361.120 176.400 ;
  LAYER ME2 ;
  RECT 1357.580 175.280 1361.120 176.400 ;
  LAYER ME1 ;
  RECT 1357.580 175.280 1361.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1348.900 175.280 1352.440 176.400 ;
  LAYER ME3 ;
  RECT 1348.900 175.280 1352.440 176.400 ;
  LAYER ME2 ;
  RECT 1348.900 175.280 1352.440 176.400 ;
  LAYER ME1 ;
  RECT 1348.900 175.280 1352.440 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1340.220 175.280 1343.760 176.400 ;
  LAYER ME3 ;
  RECT 1340.220 175.280 1343.760 176.400 ;
  LAYER ME2 ;
  RECT 1340.220 175.280 1343.760 176.400 ;
  LAYER ME1 ;
  RECT 1340.220 175.280 1343.760 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1331.540 175.280 1335.080 176.400 ;
  LAYER ME3 ;
  RECT 1331.540 175.280 1335.080 176.400 ;
  LAYER ME2 ;
  RECT 1331.540 175.280 1335.080 176.400 ;
  LAYER ME1 ;
  RECT 1331.540 175.280 1335.080 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1322.860 175.280 1326.400 176.400 ;
  LAYER ME3 ;
  RECT 1322.860 175.280 1326.400 176.400 ;
  LAYER ME2 ;
  RECT 1322.860 175.280 1326.400 176.400 ;
  LAYER ME1 ;
  RECT 1322.860 175.280 1326.400 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1314.180 175.280 1317.720 176.400 ;
  LAYER ME3 ;
  RECT 1314.180 175.280 1317.720 176.400 ;
  LAYER ME2 ;
  RECT 1314.180 175.280 1317.720 176.400 ;
  LAYER ME1 ;
  RECT 1314.180 175.280 1317.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1270.780 175.280 1274.320 176.400 ;
  LAYER ME3 ;
  RECT 1270.780 175.280 1274.320 176.400 ;
  LAYER ME2 ;
  RECT 1270.780 175.280 1274.320 176.400 ;
  LAYER ME1 ;
  RECT 1270.780 175.280 1274.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1262.100 175.280 1265.640 176.400 ;
  LAYER ME3 ;
  RECT 1262.100 175.280 1265.640 176.400 ;
  LAYER ME2 ;
  RECT 1262.100 175.280 1265.640 176.400 ;
  LAYER ME1 ;
  RECT 1262.100 175.280 1265.640 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1253.420 175.280 1256.960 176.400 ;
  LAYER ME3 ;
  RECT 1253.420 175.280 1256.960 176.400 ;
  LAYER ME2 ;
  RECT 1253.420 175.280 1256.960 176.400 ;
  LAYER ME1 ;
  RECT 1253.420 175.280 1256.960 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1244.740 175.280 1248.280 176.400 ;
  LAYER ME3 ;
  RECT 1244.740 175.280 1248.280 176.400 ;
  LAYER ME2 ;
  RECT 1244.740 175.280 1248.280 176.400 ;
  LAYER ME1 ;
  RECT 1244.740 175.280 1248.280 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1236.060 175.280 1239.600 176.400 ;
  LAYER ME3 ;
  RECT 1236.060 175.280 1239.600 176.400 ;
  LAYER ME2 ;
  RECT 1236.060 175.280 1239.600 176.400 ;
  LAYER ME1 ;
  RECT 1236.060 175.280 1239.600 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1227.380 175.280 1230.920 176.400 ;
  LAYER ME3 ;
  RECT 1227.380 175.280 1230.920 176.400 ;
  LAYER ME2 ;
  RECT 1227.380 175.280 1230.920 176.400 ;
  LAYER ME1 ;
  RECT 1227.380 175.280 1230.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1183.980 175.280 1187.520 176.400 ;
  LAYER ME3 ;
  RECT 1183.980 175.280 1187.520 176.400 ;
  LAYER ME2 ;
  RECT 1183.980 175.280 1187.520 176.400 ;
  LAYER ME1 ;
  RECT 1183.980 175.280 1187.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1175.300 175.280 1178.840 176.400 ;
  LAYER ME3 ;
  RECT 1175.300 175.280 1178.840 176.400 ;
  LAYER ME2 ;
  RECT 1175.300 175.280 1178.840 176.400 ;
  LAYER ME1 ;
  RECT 1175.300 175.280 1178.840 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1166.620 175.280 1170.160 176.400 ;
  LAYER ME3 ;
  RECT 1166.620 175.280 1170.160 176.400 ;
  LAYER ME2 ;
  RECT 1166.620 175.280 1170.160 176.400 ;
  LAYER ME1 ;
  RECT 1166.620 175.280 1170.160 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1157.940 175.280 1161.480 176.400 ;
  LAYER ME3 ;
  RECT 1157.940 175.280 1161.480 176.400 ;
  LAYER ME2 ;
  RECT 1157.940 175.280 1161.480 176.400 ;
  LAYER ME1 ;
  RECT 1157.940 175.280 1161.480 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1149.260 175.280 1152.800 176.400 ;
  LAYER ME3 ;
  RECT 1149.260 175.280 1152.800 176.400 ;
  LAYER ME2 ;
  RECT 1149.260 175.280 1152.800 176.400 ;
  LAYER ME1 ;
  RECT 1149.260 175.280 1152.800 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1140.580 175.280 1144.120 176.400 ;
  LAYER ME3 ;
  RECT 1140.580 175.280 1144.120 176.400 ;
  LAYER ME2 ;
  RECT 1140.580 175.280 1144.120 176.400 ;
  LAYER ME1 ;
  RECT 1140.580 175.280 1144.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1097.180 175.280 1100.720 176.400 ;
  LAYER ME3 ;
  RECT 1097.180 175.280 1100.720 176.400 ;
  LAYER ME2 ;
  RECT 1097.180 175.280 1100.720 176.400 ;
  LAYER ME1 ;
  RECT 1097.180 175.280 1100.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1088.500 175.280 1092.040 176.400 ;
  LAYER ME3 ;
  RECT 1088.500 175.280 1092.040 176.400 ;
  LAYER ME2 ;
  RECT 1088.500 175.280 1092.040 176.400 ;
  LAYER ME1 ;
  RECT 1088.500 175.280 1092.040 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1079.820 175.280 1083.360 176.400 ;
  LAYER ME3 ;
  RECT 1079.820 175.280 1083.360 176.400 ;
  LAYER ME2 ;
  RECT 1079.820 175.280 1083.360 176.400 ;
  LAYER ME1 ;
  RECT 1079.820 175.280 1083.360 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1071.140 175.280 1074.680 176.400 ;
  LAYER ME3 ;
  RECT 1071.140 175.280 1074.680 176.400 ;
  LAYER ME2 ;
  RECT 1071.140 175.280 1074.680 176.400 ;
  LAYER ME1 ;
  RECT 1071.140 175.280 1074.680 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1062.460 175.280 1066.000 176.400 ;
  LAYER ME3 ;
  RECT 1062.460 175.280 1066.000 176.400 ;
  LAYER ME2 ;
  RECT 1062.460 175.280 1066.000 176.400 ;
  LAYER ME1 ;
  RECT 1062.460 175.280 1066.000 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1053.780 175.280 1057.320 176.400 ;
  LAYER ME3 ;
  RECT 1053.780 175.280 1057.320 176.400 ;
  LAYER ME2 ;
  RECT 1053.780 175.280 1057.320 176.400 ;
  LAYER ME1 ;
  RECT 1053.780 175.280 1057.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1010.380 175.280 1013.920 176.400 ;
  LAYER ME3 ;
  RECT 1010.380 175.280 1013.920 176.400 ;
  LAYER ME2 ;
  RECT 1010.380 175.280 1013.920 176.400 ;
  LAYER ME1 ;
  RECT 1010.380 175.280 1013.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1001.700 175.280 1005.240 176.400 ;
  LAYER ME3 ;
  RECT 1001.700 175.280 1005.240 176.400 ;
  LAYER ME2 ;
  RECT 1001.700 175.280 1005.240 176.400 ;
  LAYER ME1 ;
  RECT 1001.700 175.280 1005.240 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.020 175.280 996.560 176.400 ;
  LAYER ME3 ;
  RECT 993.020 175.280 996.560 176.400 ;
  LAYER ME2 ;
  RECT 993.020 175.280 996.560 176.400 ;
  LAYER ME1 ;
  RECT 993.020 175.280 996.560 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 984.340 175.280 987.880 176.400 ;
  LAYER ME3 ;
  RECT 984.340 175.280 987.880 176.400 ;
  LAYER ME2 ;
  RECT 984.340 175.280 987.880 176.400 ;
  LAYER ME1 ;
  RECT 984.340 175.280 987.880 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 975.660 175.280 979.200 176.400 ;
  LAYER ME3 ;
  RECT 975.660 175.280 979.200 176.400 ;
  LAYER ME2 ;
  RECT 975.660 175.280 979.200 176.400 ;
  LAYER ME1 ;
  RECT 975.660 175.280 979.200 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 966.980 175.280 970.520 176.400 ;
  LAYER ME3 ;
  RECT 966.980 175.280 970.520 176.400 ;
  LAYER ME2 ;
  RECT 966.980 175.280 970.520 176.400 ;
  LAYER ME1 ;
  RECT 966.980 175.280 970.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 923.580 175.280 927.120 176.400 ;
  LAYER ME3 ;
  RECT 923.580 175.280 927.120 176.400 ;
  LAYER ME2 ;
  RECT 923.580 175.280 927.120 176.400 ;
  LAYER ME1 ;
  RECT 923.580 175.280 927.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 914.900 175.280 918.440 176.400 ;
  LAYER ME3 ;
  RECT 914.900 175.280 918.440 176.400 ;
  LAYER ME2 ;
  RECT 914.900 175.280 918.440 176.400 ;
  LAYER ME1 ;
  RECT 914.900 175.280 918.440 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 906.220 175.280 909.760 176.400 ;
  LAYER ME3 ;
  RECT 906.220 175.280 909.760 176.400 ;
  LAYER ME2 ;
  RECT 906.220 175.280 909.760 176.400 ;
  LAYER ME1 ;
  RECT 906.220 175.280 909.760 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 897.540 175.280 901.080 176.400 ;
  LAYER ME3 ;
  RECT 897.540 175.280 901.080 176.400 ;
  LAYER ME2 ;
  RECT 897.540 175.280 901.080 176.400 ;
  LAYER ME1 ;
  RECT 897.540 175.280 901.080 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 888.860 175.280 892.400 176.400 ;
  LAYER ME3 ;
  RECT 888.860 175.280 892.400 176.400 ;
  LAYER ME2 ;
  RECT 888.860 175.280 892.400 176.400 ;
  LAYER ME1 ;
  RECT 888.860 175.280 892.400 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 880.180 175.280 883.720 176.400 ;
  LAYER ME3 ;
  RECT 880.180 175.280 883.720 176.400 ;
  LAYER ME2 ;
  RECT 880.180 175.280 883.720 176.400 ;
  LAYER ME1 ;
  RECT 880.180 175.280 883.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 836.780 175.280 840.320 176.400 ;
  LAYER ME3 ;
  RECT 836.780 175.280 840.320 176.400 ;
  LAYER ME2 ;
  RECT 836.780 175.280 840.320 176.400 ;
  LAYER ME1 ;
  RECT 836.780 175.280 840.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 828.100 175.280 831.640 176.400 ;
  LAYER ME3 ;
  RECT 828.100 175.280 831.640 176.400 ;
  LAYER ME2 ;
  RECT 828.100 175.280 831.640 176.400 ;
  LAYER ME1 ;
  RECT 828.100 175.280 831.640 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 819.420 175.280 822.960 176.400 ;
  LAYER ME3 ;
  RECT 819.420 175.280 822.960 176.400 ;
  LAYER ME2 ;
  RECT 819.420 175.280 822.960 176.400 ;
  LAYER ME1 ;
  RECT 819.420 175.280 822.960 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 810.740 175.280 814.280 176.400 ;
  LAYER ME3 ;
  RECT 810.740 175.280 814.280 176.400 ;
  LAYER ME2 ;
  RECT 810.740 175.280 814.280 176.400 ;
  LAYER ME1 ;
  RECT 810.740 175.280 814.280 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 802.060 175.280 805.600 176.400 ;
  LAYER ME3 ;
  RECT 802.060 175.280 805.600 176.400 ;
  LAYER ME2 ;
  RECT 802.060 175.280 805.600 176.400 ;
  LAYER ME1 ;
  RECT 802.060 175.280 805.600 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 793.380 175.280 796.920 176.400 ;
  LAYER ME3 ;
  RECT 793.380 175.280 796.920 176.400 ;
  LAYER ME2 ;
  RECT 793.380 175.280 796.920 176.400 ;
  LAYER ME1 ;
  RECT 793.380 175.280 796.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 749.980 175.280 753.520 176.400 ;
  LAYER ME3 ;
  RECT 749.980 175.280 753.520 176.400 ;
  LAYER ME2 ;
  RECT 749.980 175.280 753.520 176.400 ;
  LAYER ME1 ;
  RECT 749.980 175.280 753.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 741.300 175.280 744.840 176.400 ;
  LAYER ME3 ;
  RECT 741.300 175.280 744.840 176.400 ;
  LAYER ME2 ;
  RECT 741.300 175.280 744.840 176.400 ;
  LAYER ME1 ;
  RECT 741.300 175.280 744.840 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 732.620 175.280 736.160 176.400 ;
  LAYER ME3 ;
  RECT 732.620 175.280 736.160 176.400 ;
  LAYER ME2 ;
  RECT 732.620 175.280 736.160 176.400 ;
  LAYER ME1 ;
  RECT 732.620 175.280 736.160 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 723.940 175.280 727.480 176.400 ;
  LAYER ME3 ;
  RECT 723.940 175.280 727.480 176.400 ;
  LAYER ME2 ;
  RECT 723.940 175.280 727.480 176.400 ;
  LAYER ME1 ;
  RECT 723.940 175.280 727.480 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 715.260 175.280 718.800 176.400 ;
  LAYER ME3 ;
  RECT 715.260 175.280 718.800 176.400 ;
  LAYER ME2 ;
  RECT 715.260 175.280 718.800 176.400 ;
  LAYER ME1 ;
  RECT 715.260 175.280 718.800 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 706.580 175.280 710.120 176.400 ;
  LAYER ME3 ;
  RECT 706.580 175.280 710.120 176.400 ;
  LAYER ME2 ;
  RECT 706.580 175.280 710.120 176.400 ;
  LAYER ME1 ;
  RECT 706.580 175.280 710.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 663.180 175.280 666.720 176.400 ;
  LAYER ME3 ;
  RECT 663.180 175.280 666.720 176.400 ;
  LAYER ME2 ;
  RECT 663.180 175.280 666.720 176.400 ;
  LAYER ME1 ;
  RECT 663.180 175.280 666.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.500 175.280 658.040 176.400 ;
  LAYER ME3 ;
  RECT 654.500 175.280 658.040 176.400 ;
  LAYER ME2 ;
  RECT 654.500 175.280 658.040 176.400 ;
  LAYER ME1 ;
  RECT 654.500 175.280 658.040 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 645.820 175.280 649.360 176.400 ;
  LAYER ME3 ;
  RECT 645.820 175.280 649.360 176.400 ;
  LAYER ME2 ;
  RECT 645.820 175.280 649.360 176.400 ;
  LAYER ME1 ;
  RECT 645.820 175.280 649.360 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 637.140 175.280 640.680 176.400 ;
  LAYER ME3 ;
  RECT 637.140 175.280 640.680 176.400 ;
  LAYER ME2 ;
  RECT 637.140 175.280 640.680 176.400 ;
  LAYER ME1 ;
  RECT 637.140 175.280 640.680 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 628.460 175.280 632.000 176.400 ;
  LAYER ME3 ;
  RECT 628.460 175.280 632.000 176.400 ;
  LAYER ME2 ;
  RECT 628.460 175.280 632.000 176.400 ;
  LAYER ME1 ;
  RECT 628.460 175.280 632.000 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 619.780 175.280 623.320 176.400 ;
  LAYER ME3 ;
  RECT 619.780 175.280 623.320 176.400 ;
  LAYER ME2 ;
  RECT 619.780 175.280 623.320 176.400 ;
  LAYER ME1 ;
  RECT 619.780 175.280 623.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 576.380 175.280 579.920 176.400 ;
  LAYER ME3 ;
  RECT 576.380 175.280 579.920 176.400 ;
  LAYER ME2 ;
  RECT 576.380 175.280 579.920 176.400 ;
  LAYER ME1 ;
  RECT 576.380 175.280 579.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 567.700 175.280 571.240 176.400 ;
  LAYER ME3 ;
  RECT 567.700 175.280 571.240 176.400 ;
  LAYER ME2 ;
  RECT 567.700 175.280 571.240 176.400 ;
  LAYER ME1 ;
  RECT 567.700 175.280 571.240 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 559.020 175.280 562.560 176.400 ;
  LAYER ME3 ;
  RECT 559.020 175.280 562.560 176.400 ;
  LAYER ME2 ;
  RECT 559.020 175.280 562.560 176.400 ;
  LAYER ME1 ;
  RECT 559.020 175.280 562.560 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.340 175.280 553.880 176.400 ;
  LAYER ME3 ;
  RECT 550.340 175.280 553.880 176.400 ;
  LAYER ME2 ;
  RECT 550.340 175.280 553.880 176.400 ;
  LAYER ME1 ;
  RECT 550.340 175.280 553.880 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.660 175.280 545.200 176.400 ;
  LAYER ME3 ;
  RECT 541.660 175.280 545.200 176.400 ;
  LAYER ME2 ;
  RECT 541.660 175.280 545.200 176.400 ;
  LAYER ME1 ;
  RECT 541.660 175.280 545.200 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.980 175.280 536.520 176.400 ;
  LAYER ME3 ;
  RECT 532.980 175.280 536.520 176.400 ;
  LAYER ME2 ;
  RECT 532.980 175.280 536.520 176.400 ;
  LAYER ME1 ;
  RECT 532.980 175.280 536.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.580 175.280 493.120 176.400 ;
  LAYER ME3 ;
  RECT 489.580 175.280 493.120 176.400 ;
  LAYER ME2 ;
  RECT 489.580 175.280 493.120 176.400 ;
  LAYER ME1 ;
  RECT 489.580 175.280 493.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.900 175.280 484.440 176.400 ;
  LAYER ME3 ;
  RECT 480.900 175.280 484.440 176.400 ;
  LAYER ME2 ;
  RECT 480.900 175.280 484.440 176.400 ;
  LAYER ME1 ;
  RECT 480.900 175.280 484.440 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 175.280 475.760 176.400 ;
  LAYER ME3 ;
  RECT 472.220 175.280 475.760 176.400 ;
  LAYER ME2 ;
  RECT 472.220 175.280 475.760 176.400 ;
  LAYER ME1 ;
  RECT 472.220 175.280 475.760 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.540 175.280 467.080 176.400 ;
  LAYER ME3 ;
  RECT 463.540 175.280 467.080 176.400 ;
  LAYER ME2 ;
  RECT 463.540 175.280 467.080 176.400 ;
  LAYER ME1 ;
  RECT 463.540 175.280 467.080 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.860 175.280 458.400 176.400 ;
  LAYER ME3 ;
  RECT 454.860 175.280 458.400 176.400 ;
  LAYER ME2 ;
  RECT 454.860 175.280 458.400 176.400 ;
  LAYER ME1 ;
  RECT 454.860 175.280 458.400 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.180 175.280 449.720 176.400 ;
  LAYER ME3 ;
  RECT 446.180 175.280 449.720 176.400 ;
  LAYER ME2 ;
  RECT 446.180 175.280 449.720 176.400 ;
  LAYER ME1 ;
  RECT 446.180 175.280 449.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 175.280 406.320 176.400 ;
  LAYER ME3 ;
  RECT 402.780 175.280 406.320 176.400 ;
  LAYER ME2 ;
  RECT 402.780 175.280 406.320 176.400 ;
  LAYER ME1 ;
  RECT 402.780 175.280 406.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.100 175.280 397.640 176.400 ;
  LAYER ME3 ;
  RECT 394.100 175.280 397.640 176.400 ;
  LAYER ME2 ;
  RECT 394.100 175.280 397.640 176.400 ;
  LAYER ME1 ;
  RECT 394.100 175.280 397.640 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.420 175.280 388.960 176.400 ;
  LAYER ME3 ;
  RECT 385.420 175.280 388.960 176.400 ;
  LAYER ME2 ;
  RECT 385.420 175.280 388.960 176.400 ;
  LAYER ME1 ;
  RECT 385.420 175.280 388.960 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.740 175.280 380.280 176.400 ;
  LAYER ME3 ;
  RECT 376.740 175.280 380.280 176.400 ;
  LAYER ME2 ;
  RECT 376.740 175.280 380.280 176.400 ;
  LAYER ME1 ;
  RECT 376.740 175.280 380.280 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.060 175.280 371.600 176.400 ;
  LAYER ME3 ;
  RECT 368.060 175.280 371.600 176.400 ;
  LAYER ME2 ;
  RECT 368.060 175.280 371.600 176.400 ;
  LAYER ME1 ;
  RECT 368.060 175.280 371.600 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.380 175.280 362.920 176.400 ;
  LAYER ME3 ;
  RECT 359.380 175.280 362.920 176.400 ;
  LAYER ME2 ;
  RECT 359.380 175.280 362.920 176.400 ;
  LAYER ME1 ;
  RECT 359.380 175.280 362.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.980 175.280 319.520 176.400 ;
  LAYER ME3 ;
  RECT 315.980 175.280 319.520 176.400 ;
  LAYER ME2 ;
  RECT 315.980 175.280 319.520 176.400 ;
  LAYER ME1 ;
  RECT 315.980 175.280 319.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 175.280 310.840 176.400 ;
  LAYER ME3 ;
  RECT 307.300 175.280 310.840 176.400 ;
  LAYER ME2 ;
  RECT 307.300 175.280 310.840 176.400 ;
  LAYER ME1 ;
  RECT 307.300 175.280 310.840 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 175.280 302.160 176.400 ;
  LAYER ME3 ;
  RECT 298.620 175.280 302.160 176.400 ;
  LAYER ME2 ;
  RECT 298.620 175.280 302.160 176.400 ;
  LAYER ME1 ;
  RECT 298.620 175.280 302.160 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 175.280 293.480 176.400 ;
  LAYER ME3 ;
  RECT 289.940 175.280 293.480 176.400 ;
  LAYER ME2 ;
  RECT 289.940 175.280 293.480 176.400 ;
  LAYER ME1 ;
  RECT 289.940 175.280 293.480 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 175.280 284.800 176.400 ;
  LAYER ME3 ;
  RECT 281.260 175.280 284.800 176.400 ;
  LAYER ME2 ;
  RECT 281.260 175.280 284.800 176.400 ;
  LAYER ME1 ;
  RECT 281.260 175.280 284.800 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 175.280 276.120 176.400 ;
  LAYER ME3 ;
  RECT 272.580 175.280 276.120 176.400 ;
  LAYER ME2 ;
  RECT 272.580 175.280 276.120 176.400 ;
  LAYER ME1 ;
  RECT 272.580 175.280 276.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 175.280 232.720 176.400 ;
  LAYER ME3 ;
  RECT 229.180 175.280 232.720 176.400 ;
  LAYER ME2 ;
  RECT 229.180 175.280 232.720 176.400 ;
  LAYER ME1 ;
  RECT 229.180 175.280 232.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 175.280 224.040 176.400 ;
  LAYER ME3 ;
  RECT 220.500 175.280 224.040 176.400 ;
  LAYER ME2 ;
  RECT 220.500 175.280 224.040 176.400 ;
  LAYER ME1 ;
  RECT 220.500 175.280 224.040 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 175.280 215.360 176.400 ;
  LAYER ME3 ;
  RECT 211.820 175.280 215.360 176.400 ;
  LAYER ME2 ;
  RECT 211.820 175.280 215.360 176.400 ;
  LAYER ME1 ;
  RECT 211.820 175.280 215.360 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 175.280 206.680 176.400 ;
  LAYER ME3 ;
  RECT 203.140 175.280 206.680 176.400 ;
  LAYER ME2 ;
  RECT 203.140 175.280 206.680 176.400 ;
  LAYER ME1 ;
  RECT 203.140 175.280 206.680 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 175.280 198.000 176.400 ;
  LAYER ME3 ;
  RECT 194.460 175.280 198.000 176.400 ;
  LAYER ME2 ;
  RECT 194.460 175.280 198.000 176.400 ;
  LAYER ME1 ;
  RECT 194.460 175.280 198.000 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 175.280 189.320 176.400 ;
  LAYER ME3 ;
  RECT 185.780 175.280 189.320 176.400 ;
  LAYER ME2 ;
  RECT 185.780 175.280 189.320 176.400 ;
  LAYER ME1 ;
  RECT 185.780 175.280 189.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 175.280 145.920 176.400 ;
  LAYER ME3 ;
  RECT 142.380 175.280 145.920 176.400 ;
  LAYER ME2 ;
  RECT 142.380 175.280 145.920 176.400 ;
  LAYER ME1 ;
  RECT 142.380 175.280 145.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 175.280 137.240 176.400 ;
  LAYER ME3 ;
  RECT 133.700 175.280 137.240 176.400 ;
  LAYER ME2 ;
  RECT 133.700 175.280 137.240 176.400 ;
  LAYER ME1 ;
  RECT 133.700 175.280 137.240 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 175.280 128.560 176.400 ;
  LAYER ME3 ;
  RECT 125.020 175.280 128.560 176.400 ;
  LAYER ME2 ;
  RECT 125.020 175.280 128.560 176.400 ;
  LAYER ME1 ;
  RECT 125.020 175.280 128.560 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 175.280 119.880 176.400 ;
  LAYER ME3 ;
  RECT 116.340 175.280 119.880 176.400 ;
  LAYER ME2 ;
  RECT 116.340 175.280 119.880 176.400 ;
  LAYER ME1 ;
  RECT 116.340 175.280 119.880 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 175.280 111.200 176.400 ;
  LAYER ME3 ;
  RECT 107.660 175.280 111.200 176.400 ;
  LAYER ME2 ;
  RECT 107.660 175.280 111.200 176.400 ;
  LAYER ME1 ;
  RECT 107.660 175.280 111.200 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 175.280 102.520 176.400 ;
  LAYER ME3 ;
  RECT 98.980 175.280 102.520 176.400 ;
  LAYER ME2 ;
  RECT 98.980 175.280 102.520 176.400 ;
  LAYER ME1 ;
  RECT 98.980 175.280 102.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 175.280 59.120 176.400 ;
  LAYER ME3 ;
  RECT 55.580 175.280 59.120 176.400 ;
  LAYER ME2 ;
  RECT 55.580 175.280 59.120 176.400 ;
  LAYER ME1 ;
  RECT 55.580 175.280 59.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 175.280 50.440 176.400 ;
  LAYER ME3 ;
  RECT 46.900 175.280 50.440 176.400 ;
  LAYER ME2 ;
  RECT 46.900 175.280 50.440 176.400 ;
  LAYER ME1 ;
  RECT 46.900 175.280 50.440 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 175.280 41.760 176.400 ;
  LAYER ME3 ;
  RECT 38.220 175.280 41.760 176.400 ;
  LAYER ME2 ;
  RECT 38.220 175.280 41.760 176.400 ;
  LAYER ME1 ;
  RECT 38.220 175.280 41.760 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 175.280 33.080 176.400 ;
  LAYER ME3 ;
  RECT 29.540 175.280 33.080 176.400 ;
  LAYER ME2 ;
  RECT 29.540 175.280 33.080 176.400 ;
  LAYER ME1 ;
  RECT 29.540 175.280 33.080 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 175.280 24.400 176.400 ;
  LAYER ME3 ;
  RECT 20.860 175.280 24.400 176.400 ;
  LAYER ME2 ;
  RECT 20.860 175.280 24.400 176.400 ;
  LAYER ME1 ;
  RECT 20.860 175.280 24.400 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 175.280 15.720 176.400 ;
  LAYER ME3 ;
  RECT 12.180 175.280 15.720 176.400 ;
  LAYER ME2 ;
  RECT 12.180 175.280 15.720 176.400 ;
  LAYER ME1 ;
  RECT 12.180 175.280 15.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1879.000 0.000 1882.540 1.120 ;
  LAYER ME3 ;
  RECT 1879.000 0.000 1882.540 1.120 ;
  LAYER ME2 ;
  RECT 1879.000 0.000 1882.540 1.120 ;
  LAYER ME1 ;
  RECT 1879.000 0.000 1882.540 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1857.300 0.000 1860.840 1.120 ;
  LAYER ME3 ;
  RECT 1857.300 0.000 1860.840 1.120 ;
  LAYER ME2 ;
  RECT 1857.300 0.000 1860.840 1.120 ;
  LAYER ME1 ;
  RECT 1857.300 0.000 1860.840 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1835.600 0.000 1839.140 1.120 ;
  LAYER ME3 ;
  RECT 1835.600 0.000 1839.140 1.120 ;
  LAYER ME2 ;
  RECT 1835.600 0.000 1839.140 1.120 ;
  LAYER ME1 ;
  RECT 1835.600 0.000 1839.140 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1809.560 0.000 1813.100 1.120 ;
  LAYER ME3 ;
  RECT 1809.560 0.000 1813.100 1.120 ;
  LAYER ME2 ;
  RECT 1809.560 0.000 1813.100 1.120 ;
  LAYER ME1 ;
  RECT 1809.560 0.000 1813.100 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1696.100 0.000 1699.640 1.120 ;
  LAYER ME3 ;
  RECT 1696.100 0.000 1699.640 1.120 ;
  LAYER ME2 ;
  RECT 1696.100 0.000 1699.640 1.120 ;
  LAYER ME1 ;
  RECT 1696.100 0.000 1699.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1679.360 0.000 1682.900 1.120 ;
  LAYER ME3 ;
  RECT 1679.360 0.000 1682.900 1.120 ;
  LAYER ME2 ;
  RECT 1679.360 0.000 1682.900 1.120 ;
  LAYER ME1 ;
  RECT 1679.360 0.000 1682.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1652.700 0.000 1656.240 1.120 ;
  LAYER ME3 ;
  RECT 1652.700 0.000 1656.240 1.120 ;
  LAYER ME2 ;
  RECT 1652.700 0.000 1656.240 1.120 ;
  LAYER ME1 ;
  RECT 1652.700 0.000 1656.240 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1631.620 0.000 1635.160 1.120 ;
  LAYER ME3 ;
  RECT 1631.620 0.000 1635.160 1.120 ;
  LAYER ME2 ;
  RECT 1631.620 0.000 1635.160 1.120 ;
  LAYER ME1 ;
  RECT 1631.620 0.000 1635.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1609.920 0.000 1613.460 1.120 ;
  LAYER ME3 ;
  RECT 1609.920 0.000 1613.460 1.120 ;
  LAYER ME2 ;
  RECT 1609.920 0.000 1613.460 1.120 ;
  LAYER ME1 ;
  RECT 1609.920 0.000 1613.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1583.260 0.000 1586.800 1.120 ;
  LAYER ME3 ;
  RECT 1583.260 0.000 1586.800 1.120 ;
  LAYER ME2 ;
  RECT 1583.260 0.000 1586.800 1.120 ;
  LAYER ME1 ;
  RECT 1583.260 0.000 1586.800 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1470.420 0.000 1473.960 1.120 ;
  LAYER ME3 ;
  RECT 1470.420 0.000 1473.960 1.120 ;
  LAYER ME2 ;
  RECT 1470.420 0.000 1473.960 1.120 ;
  LAYER ME1 ;
  RECT 1470.420 0.000 1473.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1453.680 0.000 1457.220 1.120 ;
  LAYER ME3 ;
  RECT 1453.680 0.000 1457.220 1.120 ;
  LAYER ME2 ;
  RECT 1453.680 0.000 1457.220 1.120 ;
  LAYER ME1 ;
  RECT 1453.680 0.000 1457.220 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1427.020 0.000 1430.560 1.120 ;
  LAYER ME3 ;
  RECT 1427.020 0.000 1430.560 1.120 ;
  LAYER ME2 ;
  RECT 1427.020 0.000 1430.560 1.120 ;
  LAYER ME1 ;
  RECT 1427.020 0.000 1430.560 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1405.320 0.000 1408.860 1.120 ;
  LAYER ME3 ;
  RECT 1405.320 0.000 1408.860 1.120 ;
  LAYER ME2 ;
  RECT 1405.320 0.000 1408.860 1.120 ;
  LAYER ME1 ;
  RECT 1405.320 0.000 1408.860 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1383.620 0.000 1387.160 1.120 ;
  LAYER ME3 ;
  RECT 1383.620 0.000 1387.160 1.120 ;
  LAYER ME2 ;
  RECT 1383.620 0.000 1387.160 1.120 ;
  LAYER ME1 ;
  RECT 1383.620 0.000 1387.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1356.960 0.000 1360.500 1.120 ;
  LAYER ME3 ;
  RECT 1356.960 0.000 1360.500 1.120 ;
  LAYER ME2 ;
  RECT 1356.960 0.000 1360.500 1.120 ;
  LAYER ME1 ;
  RECT 1356.960 0.000 1360.500 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1244.120 0.000 1247.660 1.120 ;
  LAYER ME3 ;
  RECT 1244.120 0.000 1247.660 1.120 ;
  LAYER ME2 ;
  RECT 1244.120 0.000 1247.660 1.120 ;
  LAYER ME1 ;
  RECT 1244.120 0.000 1247.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1227.380 0.000 1230.920 1.120 ;
  LAYER ME3 ;
  RECT 1227.380 0.000 1230.920 1.120 ;
  LAYER ME2 ;
  RECT 1227.380 0.000 1230.920 1.120 ;
  LAYER ME1 ;
  RECT 1227.380 0.000 1230.920 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1200.720 0.000 1204.260 1.120 ;
  LAYER ME3 ;
  RECT 1200.720 0.000 1204.260 1.120 ;
  LAYER ME2 ;
  RECT 1200.720 0.000 1204.260 1.120 ;
  LAYER ME1 ;
  RECT 1200.720 0.000 1204.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1179.020 0.000 1182.560 1.120 ;
  LAYER ME3 ;
  RECT 1179.020 0.000 1182.560 1.120 ;
  LAYER ME2 ;
  RECT 1179.020 0.000 1182.560 1.120 ;
  LAYER ME1 ;
  RECT 1179.020 0.000 1182.560 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER ME3 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER ME2 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER ME1 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1131.280 0.000 1134.820 1.120 ;
  LAYER ME3 ;
  RECT 1131.280 0.000 1134.820 1.120 ;
  LAYER ME2 ;
  RECT 1131.280 0.000 1134.820 1.120 ;
  LAYER ME1 ;
  RECT 1131.280 0.000 1134.820 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1017.820 0.000 1021.360 1.120 ;
  LAYER ME3 ;
  RECT 1017.820 0.000 1021.360 1.120 ;
  LAYER ME2 ;
  RECT 1017.820 0.000 1021.360 1.120 ;
  LAYER ME1 ;
  RECT 1017.820 0.000 1021.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1001.080 0.000 1004.620 1.120 ;
  LAYER ME3 ;
  RECT 1001.080 0.000 1004.620 1.120 ;
  LAYER ME2 ;
  RECT 1001.080 0.000 1004.620 1.120 ;
  LAYER ME1 ;
  RECT 1001.080 0.000 1004.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER ME3 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER ME2 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER ME1 ;
  RECT 965.120 0.000 968.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER ME3 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER ME2 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER ME1 ;
  RECT 956.440 0.000 959.980 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 935.360 0.000 938.900 1.120 ;
  LAYER ME3 ;
  RECT 935.360 0.000 938.900 1.120 ;
  LAYER ME2 ;
  RECT 935.360 0.000 938.900 1.120 ;
  LAYER ME1 ;
  RECT 935.360 0.000 938.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 917.380 0.000 920.920 1.120 ;
  LAYER ME3 ;
  RECT 917.380 0.000 920.920 1.120 ;
  LAYER ME2 ;
  RECT 917.380 0.000 920.920 1.120 ;
  LAYER ME1 ;
  RECT 917.380 0.000 920.920 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 818.180 0.000 821.720 1.120 ;
  LAYER ME3 ;
  RECT 818.180 0.000 821.720 1.120 ;
  LAYER ME2 ;
  RECT 818.180 0.000 821.720 1.120 ;
  LAYER ME1 ;
  RECT 818.180 0.000 821.720 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 792.140 0.000 795.680 1.120 ;
  LAYER ME3 ;
  RECT 792.140 0.000 795.680 1.120 ;
  LAYER ME2 ;
  RECT 792.140 0.000 795.680 1.120 ;
  LAYER ME1 ;
  RECT 792.140 0.000 795.680 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER ME3 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER ME2 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER ME1 ;
  RECT 770.440 0.000 773.980 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER ME3 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER ME2 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER ME1 ;
  RECT 748.740 0.000 752.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 722.080 0.000 725.620 1.120 ;
  LAYER ME3 ;
  RECT 722.080 0.000 725.620 1.120 ;
  LAYER ME2 ;
  RECT 722.080 0.000 725.620 1.120 ;
  LAYER ME1 ;
  RECT 722.080 0.000 725.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 705.340 0.000 708.880 1.120 ;
  LAYER ME3 ;
  RECT 705.340 0.000 708.880 1.120 ;
  LAYER ME2 ;
  RECT 705.340 0.000 708.880 1.120 ;
  LAYER ME1 ;
  RECT 705.340 0.000 708.880 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER ME3 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER ME2 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER ME1 ;
  RECT 592.500 0.000 596.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER ME3 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER ME2 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER ME1 ;
  RECT 544.140 0.000 547.680 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME3 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME2 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME1 ;
  RECT 522.440 0.000 525.980 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.780 0.000 499.320 1.120 ;
  LAYER ME3 ;
  RECT 495.780 0.000 499.320 1.120 ;
  LAYER ME2 ;
  RECT 495.780 0.000 499.320 1.120 ;
  LAYER ME1 ;
  RECT 495.780 0.000 499.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER ME3 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER ME2 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER ME1 ;
  RECT 479.040 0.000 482.580 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER ME3 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER ME2 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER ME1 ;
  RECT 366.200 0.000 369.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME3 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME2 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME1 ;
  RECT 318.460 0.000 322.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME3 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME2 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME1 ;
  RECT 296.760 0.000 300.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME3 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME2 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME1 ;
  RECT 270.100 0.000 273.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO127
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1885.480 0.000 1886.600 1.120 ;
  LAYER ME3 ;
  RECT 1885.480 0.000 1886.600 1.120 ;
  LAYER ME2 ;
  RECT 1885.480 0.000 1886.600 1.120 ;
  LAYER ME1 ;
  RECT 1885.480 0.000 1886.600 1.120 ;
 END
END DO127
PIN DI127
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1876.800 0.000 1877.920 1.120 ;
  LAYER ME3 ;
  RECT 1876.800 0.000 1877.920 1.120 ;
  LAYER ME2 ;
  RECT 1876.800 0.000 1877.920 1.120 ;
  LAYER ME1 ;
  RECT 1876.800 0.000 1877.920 1.120 ;
 END
END DI127
PIN DO126
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1871.840 0.000 1872.960 1.120 ;
  LAYER ME3 ;
  RECT 1871.840 0.000 1872.960 1.120 ;
  LAYER ME2 ;
  RECT 1871.840 0.000 1872.960 1.120 ;
  LAYER ME1 ;
  RECT 1871.840 0.000 1872.960 1.120 ;
 END
END DO126
PIN DI126
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1863.780 0.000 1864.900 1.120 ;
  LAYER ME3 ;
  RECT 1863.780 0.000 1864.900 1.120 ;
  LAYER ME2 ;
  RECT 1863.780 0.000 1864.900 1.120 ;
  LAYER ME1 ;
  RECT 1863.780 0.000 1864.900 1.120 ;
 END
END DI126
PIN DO125
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1855.100 0.000 1856.220 1.120 ;
  LAYER ME3 ;
  RECT 1855.100 0.000 1856.220 1.120 ;
  LAYER ME2 ;
  RECT 1855.100 0.000 1856.220 1.120 ;
  LAYER ME1 ;
  RECT 1855.100 0.000 1856.220 1.120 ;
 END
END DO125
PIN DI125
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1847.040 0.000 1848.160 1.120 ;
  LAYER ME3 ;
  RECT 1847.040 0.000 1848.160 1.120 ;
  LAYER ME2 ;
  RECT 1847.040 0.000 1848.160 1.120 ;
  LAYER ME1 ;
  RECT 1847.040 0.000 1848.160 1.120 ;
 END
END DI125
PIN DO124
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER ME3 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER ME2 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER ME1 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
 END
END DO124
PIN DI124
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
  LAYER ME3 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
  LAYER ME2 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
  LAYER ME1 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
 END
END DI124
PIN DO123
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1829.060 0.000 1830.180 1.120 ;
  LAYER ME3 ;
  RECT 1829.060 0.000 1830.180 1.120 ;
  LAYER ME2 ;
  RECT 1829.060 0.000 1830.180 1.120 ;
  LAYER ME1 ;
  RECT 1829.060 0.000 1830.180 1.120 ;
 END
END DO123
PIN DI123
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1820.380 0.000 1821.500 1.120 ;
  LAYER ME3 ;
  RECT 1820.380 0.000 1821.500 1.120 ;
  LAYER ME2 ;
  RECT 1820.380 0.000 1821.500 1.120 ;
  LAYER ME1 ;
  RECT 1820.380 0.000 1821.500 1.120 ;
 END
END DI123
PIN DO122
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
  LAYER ME3 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
  LAYER ME2 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
  LAYER ME1 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
 END
END DO122
PIN DI122
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1807.360 0.000 1808.480 1.120 ;
  LAYER ME3 ;
  RECT 1807.360 0.000 1808.480 1.120 ;
  LAYER ME2 ;
  RECT 1807.360 0.000 1808.480 1.120 ;
  LAYER ME1 ;
  RECT 1807.360 0.000 1808.480 1.120 ;
 END
END DI122
PIN DO121
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1798.680 0.000 1799.800 1.120 ;
  LAYER ME3 ;
  RECT 1798.680 0.000 1799.800 1.120 ;
  LAYER ME2 ;
  RECT 1798.680 0.000 1799.800 1.120 ;
  LAYER ME1 ;
  RECT 1798.680 0.000 1799.800 1.120 ;
 END
END DO121
PIN DI121
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER ME3 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER ME2 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER ME1 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
 END
END DI121
PIN DO120
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1785.660 0.000 1786.780 1.120 ;
  LAYER ME3 ;
  RECT 1785.660 0.000 1786.780 1.120 ;
  LAYER ME2 ;
  RECT 1785.660 0.000 1786.780 1.120 ;
  LAYER ME1 ;
  RECT 1785.660 0.000 1786.780 1.120 ;
 END
END DO120
PIN DI120
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1776.980 0.000 1778.100 1.120 ;
  LAYER ME3 ;
  RECT 1776.980 0.000 1778.100 1.120 ;
  LAYER ME2 ;
  RECT 1776.980 0.000 1778.100 1.120 ;
  LAYER ME1 ;
  RECT 1776.980 0.000 1778.100 1.120 ;
 END
END DI120
PIN DO119
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER ME3 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER ME2 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER ME1 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
 END
END DO119
PIN DI119
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
  LAYER ME3 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
  LAYER ME2 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
  LAYER ME1 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
 END
END DI119
PIN DO118
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1759.000 0.000 1760.120 1.120 ;
  LAYER ME3 ;
  RECT 1759.000 0.000 1760.120 1.120 ;
  LAYER ME2 ;
  RECT 1759.000 0.000 1760.120 1.120 ;
  LAYER ME1 ;
  RECT 1759.000 0.000 1760.120 1.120 ;
 END
END DO118
PIN DI118
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1750.320 0.000 1751.440 1.120 ;
  LAYER ME3 ;
  RECT 1750.320 0.000 1751.440 1.120 ;
  LAYER ME2 ;
  RECT 1750.320 0.000 1751.440 1.120 ;
  LAYER ME1 ;
  RECT 1750.320 0.000 1751.440 1.120 ;
 END
END DI118
PIN DO117
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1742.260 0.000 1743.380 1.120 ;
  LAYER ME3 ;
  RECT 1742.260 0.000 1743.380 1.120 ;
  LAYER ME2 ;
  RECT 1742.260 0.000 1743.380 1.120 ;
  LAYER ME1 ;
  RECT 1742.260 0.000 1743.380 1.120 ;
 END
END DO117
PIN DI117
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1733.580 0.000 1734.700 1.120 ;
  LAYER ME3 ;
  RECT 1733.580 0.000 1734.700 1.120 ;
  LAYER ME2 ;
  RECT 1733.580 0.000 1734.700 1.120 ;
  LAYER ME1 ;
  RECT 1733.580 0.000 1734.700 1.120 ;
 END
END DI117
PIN DO116
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1729.240 0.000 1730.360 1.120 ;
  LAYER ME3 ;
  RECT 1729.240 0.000 1730.360 1.120 ;
  LAYER ME2 ;
  RECT 1729.240 0.000 1730.360 1.120 ;
  LAYER ME1 ;
  RECT 1729.240 0.000 1730.360 1.120 ;
 END
END DO116
PIN DI116
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1720.560 0.000 1721.680 1.120 ;
  LAYER ME3 ;
  RECT 1720.560 0.000 1721.680 1.120 ;
  LAYER ME2 ;
  RECT 1720.560 0.000 1721.680 1.120 ;
  LAYER ME1 ;
  RECT 1720.560 0.000 1721.680 1.120 ;
 END
END DI116
PIN DO115
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1715.600 0.000 1716.720 1.120 ;
  LAYER ME3 ;
  RECT 1715.600 0.000 1716.720 1.120 ;
  LAYER ME2 ;
  RECT 1715.600 0.000 1716.720 1.120 ;
  LAYER ME1 ;
  RECT 1715.600 0.000 1716.720 1.120 ;
 END
END DO115
PIN DI115
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1707.540 0.000 1708.660 1.120 ;
  LAYER ME3 ;
  RECT 1707.540 0.000 1708.660 1.120 ;
  LAYER ME2 ;
  RECT 1707.540 0.000 1708.660 1.120 ;
  LAYER ME1 ;
  RECT 1707.540 0.000 1708.660 1.120 ;
 END
END DI115
PIN DO114
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1702.580 0.000 1703.700 1.120 ;
  LAYER ME3 ;
  RECT 1702.580 0.000 1703.700 1.120 ;
  LAYER ME2 ;
  RECT 1702.580 0.000 1703.700 1.120 ;
  LAYER ME1 ;
  RECT 1702.580 0.000 1703.700 1.120 ;
 END
END DO114
PIN DI114
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1693.900 0.000 1695.020 1.120 ;
  LAYER ME3 ;
  RECT 1693.900 0.000 1695.020 1.120 ;
  LAYER ME2 ;
  RECT 1693.900 0.000 1695.020 1.120 ;
  LAYER ME1 ;
  RECT 1693.900 0.000 1695.020 1.120 ;
 END
END DI114
PIN DO113
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1685.840 0.000 1686.960 1.120 ;
  LAYER ME3 ;
  RECT 1685.840 0.000 1686.960 1.120 ;
  LAYER ME2 ;
  RECT 1685.840 0.000 1686.960 1.120 ;
  LAYER ME1 ;
  RECT 1685.840 0.000 1686.960 1.120 ;
 END
END DO113
PIN DI113
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1677.160 0.000 1678.280 1.120 ;
  LAYER ME3 ;
  RECT 1677.160 0.000 1678.280 1.120 ;
  LAYER ME2 ;
  RECT 1677.160 0.000 1678.280 1.120 ;
  LAYER ME1 ;
  RECT 1677.160 0.000 1678.280 1.120 ;
 END
END DI113
PIN DO112
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1672.200 0.000 1673.320 1.120 ;
  LAYER ME3 ;
  RECT 1672.200 0.000 1673.320 1.120 ;
  LAYER ME2 ;
  RECT 1672.200 0.000 1673.320 1.120 ;
  LAYER ME1 ;
  RECT 1672.200 0.000 1673.320 1.120 ;
 END
END DO112
PIN DI112
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1664.140 0.000 1665.260 1.120 ;
  LAYER ME3 ;
  RECT 1664.140 0.000 1665.260 1.120 ;
  LAYER ME2 ;
  RECT 1664.140 0.000 1665.260 1.120 ;
  LAYER ME1 ;
  RECT 1664.140 0.000 1665.260 1.120 ;
 END
END DI112
PIN DO111
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1659.180 0.000 1660.300 1.120 ;
  LAYER ME3 ;
  RECT 1659.180 0.000 1660.300 1.120 ;
  LAYER ME2 ;
  RECT 1659.180 0.000 1660.300 1.120 ;
  LAYER ME1 ;
  RECT 1659.180 0.000 1660.300 1.120 ;
 END
END DO111
PIN DI111
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1650.500 0.000 1651.620 1.120 ;
  LAYER ME3 ;
  RECT 1650.500 0.000 1651.620 1.120 ;
  LAYER ME2 ;
  RECT 1650.500 0.000 1651.620 1.120 ;
  LAYER ME1 ;
  RECT 1650.500 0.000 1651.620 1.120 ;
 END
END DI111
PIN DO110
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1646.160 0.000 1647.280 1.120 ;
  LAYER ME3 ;
  RECT 1646.160 0.000 1647.280 1.120 ;
  LAYER ME2 ;
  RECT 1646.160 0.000 1647.280 1.120 ;
  LAYER ME1 ;
  RECT 1646.160 0.000 1647.280 1.120 ;
 END
END DO110
PIN DI110
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1637.480 0.000 1638.600 1.120 ;
  LAYER ME3 ;
  RECT 1637.480 0.000 1638.600 1.120 ;
  LAYER ME2 ;
  RECT 1637.480 0.000 1638.600 1.120 ;
  LAYER ME1 ;
  RECT 1637.480 0.000 1638.600 1.120 ;
 END
END DI110
PIN DO109
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1629.420 0.000 1630.540 1.120 ;
  LAYER ME3 ;
  RECT 1629.420 0.000 1630.540 1.120 ;
  LAYER ME2 ;
  RECT 1629.420 0.000 1630.540 1.120 ;
  LAYER ME1 ;
  RECT 1629.420 0.000 1630.540 1.120 ;
 END
END DO109
PIN DI109
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1620.740 0.000 1621.860 1.120 ;
  LAYER ME3 ;
  RECT 1620.740 0.000 1621.860 1.120 ;
  LAYER ME2 ;
  RECT 1620.740 0.000 1621.860 1.120 ;
  LAYER ME1 ;
  RECT 1620.740 0.000 1621.860 1.120 ;
 END
END DI109
PIN DO108
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1615.780 0.000 1616.900 1.120 ;
  LAYER ME3 ;
  RECT 1615.780 0.000 1616.900 1.120 ;
  LAYER ME2 ;
  RECT 1615.780 0.000 1616.900 1.120 ;
  LAYER ME1 ;
  RECT 1615.780 0.000 1616.900 1.120 ;
 END
END DO108
PIN DI108
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1607.720 0.000 1608.840 1.120 ;
  LAYER ME3 ;
  RECT 1607.720 0.000 1608.840 1.120 ;
  LAYER ME2 ;
  RECT 1607.720 0.000 1608.840 1.120 ;
  LAYER ME1 ;
  RECT 1607.720 0.000 1608.840 1.120 ;
 END
END DI108
PIN DO107
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1602.760 0.000 1603.880 1.120 ;
  LAYER ME3 ;
  RECT 1602.760 0.000 1603.880 1.120 ;
  LAYER ME2 ;
  RECT 1602.760 0.000 1603.880 1.120 ;
  LAYER ME1 ;
  RECT 1602.760 0.000 1603.880 1.120 ;
 END
END DO107
PIN DI107
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1594.080 0.000 1595.200 1.120 ;
  LAYER ME3 ;
  RECT 1594.080 0.000 1595.200 1.120 ;
  LAYER ME2 ;
  RECT 1594.080 0.000 1595.200 1.120 ;
  LAYER ME1 ;
  RECT 1594.080 0.000 1595.200 1.120 ;
 END
END DI107
PIN DO106
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1589.120 0.000 1590.240 1.120 ;
  LAYER ME3 ;
  RECT 1589.120 0.000 1590.240 1.120 ;
  LAYER ME2 ;
  RECT 1589.120 0.000 1590.240 1.120 ;
  LAYER ME1 ;
  RECT 1589.120 0.000 1590.240 1.120 ;
 END
END DO106
PIN DI106
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1581.060 0.000 1582.180 1.120 ;
  LAYER ME3 ;
  RECT 1581.060 0.000 1582.180 1.120 ;
  LAYER ME2 ;
  RECT 1581.060 0.000 1582.180 1.120 ;
  LAYER ME1 ;
  RECT 1581.060 0.000 1582.180 1.120 ;
 END
END DI106
PIN DO105
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1573.000 0.000 1574.120 1.120 ;
  LAYER ME3 ;
  RECT 1573.000 0.000 1574.120 1.120 ;
  LAYER ME2 ;
  RECT 1573.000 0.000 1574.120 1.120 ;
  LAYER ME1 ;
  RECT 1573.000 0.000 1574.120 1.120 ;
 END
END DO105
PIN DI105
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1564.320 0.000 1565.440 1.120 ;
  LAYER ME3 ;
  RECT 1564.320 0.000 1565.440 1.120 ;
  LAYER ME2 ;
  RECT 1564.320 0.000 1565.440 1.120 ;
  LAYER ME1 ;
  RECT 1564.320 0.000 1565.440 1.120 ;
 END
END DI105
PIN DO104
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1559.360 0.000 1560.480 1.120 ;
  LAYER ME3 ;
  RECT 1559.360 0.000 1560.480 1.120 ;
  LAYER ME2 ;
  RECT 1559.360 0.000 1560.480 1.120 ;
  LAYER ME1 ;
  RECT 1559.360 0.000 1560.480 1.120 ;
 END
END DO104
PIN DI104
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1551.300 0.000 1552.420 1.120 ;
  LAYER ME3 ;
  RECT 1551.300 0.000 1552.420 1.120 ;
  LAYER ME2 ;
  RECT 1551.300 0.000 1552.420 1.120 ;
  LAYER ME1 ;
  RECT 1551.300 0.000 1552.420 1.120 ;
 END
END DI104
PIN DO103
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1546.340 0.000 1547.460 1.120 ;
  LAYER ME3 ;
  RECT 1546.340 0.000 1547.460 1.120 ;
  LAYER ME2 ;
  RECT 1546.340 0.000 1547.460 1.120 ;
  LAYER ME1 ;
  RECT 1546.340 0.000 1547.460 1.120 ;
 END
END DO103
PIN DI103
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1537.660 0.000 1538.780 1.120 ;
  LAYER ME3 ;
  RECT 1537.660 0.000 1538.780 1.120 ;
  LAYER ME2 ;
  RECT 1537.660 0.000 1538.780 1.120 ;
  LAYER ME1 ;
  RECT 1537.660 0.000 1538.780 1.120 ;
 END
END DI103
PIN DO102
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1532.700 0.000 1533.820 1.120 ;
  LAYER ME3 ;
  RECT 1532.700 0.000 1533.820 1.120 ;
  LAYER ME2 ;
  RECT 1532.700 0.000 1533.820 1.120 ;
  LAYER ME1 ;
  RECT 1532.700 0.000 1533.820 1.120 ;
 END
END DO102
PIN DI102
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1524.640 0.000 1525.760 1.120 ;
  LAYER ME3 ;
  RECT 1524.640 0.000 1525.760 1.120 ;
  LAYER ME2 ;
  RECT 1524.640 0.000 1525.760 1.120 ;
  LAYER ME1 ;
  RECT 1524.640 0.000 1525.760 1.120 ;
 END
END DI102
PIN DO101
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1515.960 0.000 1517.080 1.120 ;
  LAYER ME3 ;
  RECT 1515.960 0.000 1517.080 1.120 ;
  LAYER ME2 ;
  RECT 1515.960 0.000 1517.080 1.120 ;
  LAYER ME1 ;
  RECT 1515.960 0.000 1517.080 1.120 ;
 END
END DO101
PIN DI101
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1507.900 0.000 1509.020 1.120 ;
  LAYER ME3 ;
  RECT 1507.900 0.000 1509.020 1.120 ;
  LAYER ME2 ;
  RECT 1507.900 0.000 1509.020 1.120 ;
  LAYER ME1 ;
  RECT 1507.900 0.000 1509.020 1.120 ;
 END
END DI101
PIN DO100
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1502.940 0.000 1504.060 1.120 ;
  LAYER ME3 ;
  RECT 1502.940 0.000 1504.060 1.120 ;
  LAYER ME2 ;
  RECT 1502.940 0.000 1504.060 1.120 ;
  LAYER ME1 ;
  RECT 1502.940 0.000 1504.060 1.120 ;
 END
END DO100
PIN DI100
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1494.260 0.000 1495.380 1.120 ;
  LAYER ME3 ;
  RECT 1494.260 0.000 1495.380 1.120 ;
  LAYER ME2 ;
  RECT 1494.260 0.000 1495.380 1.120 ;
  LAYER ME1 ;
  RECT 1494.260 0.000 1495.380 1.120 ;
 END
END DI100
PIN DO99
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1489.920 0.000 1491.040 1.120 ;
  LAYER ME3 ;
  RECT 1489.920 0.000 1491.040 1.120 ;
  LAYER ME2 ;
  RECT 1489.920 0.000 1491.040 1.120 ;
  LAYER ME1 ;
  RECT 1489.920 0.000 1491.040 1.120 ;
 END
END DO99
PIN DI99
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1481.240 0.000 1482.360 1.120 ;
  LAYER ME3 ;
  RECT 1481.240 0.000 1482.360 1.120 ;
  LAYER ME2 ;
  RECT 1481.240 0.000 1482.360 1.120 ;
  LAYER ME1 ;
  RECT 1481.240 0.000 1482.360 1.120 ;
 END
END DI99
PIN DO98
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1476.280 0.000 1477.400 1.120 ;
  LAYER ME3 ;
  RECT 1476.280 0.000 1477.400 1.120 ;
  LAYER ME2 ;
  RECT 1476.280 0.000 1477.400 1.120 ;
  LAYER ME1 ;
  RECT 1476.280 0.000 1477.400 1.120 ;
 END
END DO98
PIN DI98
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1468.220 0.000 1469.340 1.120 ;
  LAYER ME3 ;
  RECT 1468.220 0.000 1469.340 1.120 ;
  LAYER ME2 ;
  RECT 1468.220 0.000 1469.340 1.120 ;
  LAYER ME1 ;
  RECT 1468.220 0.000 1469.340 1.120 ;
 END
END DI98
PIN DO97
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1459.540 0.000 1460.660 1.120 ;
  LAYER ME3 ;
  RECT 1459.540 0.000 1460.660 1.120 ;
  LAYER ME2 ;
  RECT 1459.540 0.000 1460.660 1.120 ;
  LAYER ME1 ;
  RECT 1459.540 0.000 1460.660 1.120 ;
 END
END DO97
PIN DI97
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1451.480 0.000 1452.600 1.120 ;
  LAYER ME3 ;
  RECT 1451.480 0.000 1452.600 1.120 ;
  LAYER ME2 ;
  RECT 1451.480 0.000 1452.600 1.120 ;
  LAYER ME1 ;
  RECT 1451.480 0.000 1452.600 1.120 ;
 END
END DI97
PIN DO96
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1446.520 0.000 1447.640 1.120 ;
  LAYER ME3 ;
  RECT 1446.520 0.000 1447.640 1.120 ;
  LAYER ME2 ;
  RECT 1446.520 0.000 1447.640 1.120 ;
  LAYER ME1 ;
  RECT 1446.520 0.000 1447.640 1.120 ;
 END
END DO96
PIN DI96
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1437.840 0.000 1438.960 1.120 ;
  LAYER ME3 ;
  RECT 1437.840 0.000 1438.960 1.120 ;
  LAYER ME2 ;
  RECT 1437.840 0.000 1438.960 1.120 ;
  LAYER ME1 ;
  RECT 1437.840 0.000 1438.960 1.120 ;
 END
END DI96
PIN DO95
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1432.880 0.000 1434.000 1.120 ;
  LAYER ME3 ;
  RECT 1432.880 0.000 1434.000 1.120 ;
  LAYER ME2 ;
  RECT 1432.880 0.000 1434.000 1.120 ;
  LAYER ME1 ;
  RECT 1432.880 0.000 1434.000 1.120 ;
 END
END DO95
PIN DI95
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1424.820 0.000 1425.940 1.120 ;
  LAYER ME3 ;
  RECT 1424.820 0.000 1425.940 1.120 ;
  LAYER ME2 ;
  RECT 1424.820 0.000 1425.940 1.120 ;
  LAYER ME1 ;
  RECT 1424.820 0.000 1425.940 1.120 ;
 END
END DI95
PIN DO94
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1419.860 0.000 1420.980 1.120 ;
  LAYER ME3 ;
  RECT 1419.860 0.000 1420.980 1.120 ;
  LAYER ME2 ;
  RECT 1419.860 0.000 1420.980 1.120 ;
  LAYER ME1 ;
  RECT 1419.860 0.000 1420.980 1.120 ;
 END
END DO94
PIN DI94
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1411.180 0.000 1412.300 1.120 ;
  LAYER ME3 ;
  RECT 1411.180 0.000 1412.300 1.120 ;
  LAYER ME2 ;
  RECT 1411.180 0.000 1412.300 1.120 ;
  LAYER ME1 ;
  RECT 1411.180 0.000 1412.300 1.120 ;
 END
END DI94
PIN DO93
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1403.120 0.000 1404.240 1.120 ;
  LAYER ME3 ;
  RECT 1403.120 0.000 1404.240 1.120 ;
  LAYER ME2 ;
  RECT 1403.120 0.000 1404.240 1.120 ;
  LAYER ME1 ;
  RECT 1403.120 0.000 1404.240 1.120 ;
 END
END DO93
PIN DI93
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1395.060 0.000 1396.180 1.120 ;
  LAYER ME3 ;
  RECT 1395.060 0.000 1396.180 1.120 ;
  LAYER ME2 ;
  RECT 1395.060 0.000 1396.180 1.120 ;
  LAYER ME1 ;
  RECT 1395.060 0.000 1396.180 1.120 ;
 END
END DI93
PIN DO92
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1390.100 0.000 1391.220 1.120 ;
  LAYER ME3 ;
  RECT 1390.100 0.000 1391.220 1.120 ;
  LAYER ME2 ;
  RECT 1390.100 0.000 1391.220 1.120 ;
  LAYER ME1 ;
  RECT 1390.100 0.000 1391.220 1.120 ;
 END
END DO92
PIN DI92
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1381.420 0.000 1382.540 1.120 ;
  LAYER ME3 ;
  RECT 1381.420 0.000 1382.540 1.120 ;
  LAYER ME2 ;
  RECT 1381.420 0.000 1382.540 1.120 ;
  LAYER ME1 ;
  RECT 1381.420 0.000 1382.540 1.120 ;
 END
END DI92
PIN DO91
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1376.460 0.000 1377.580 1.120 ;
  LAYER ME3 ;
  RECT 1376.460 0.000 1377.580 1.120 ;
  LAYER ME2 ;
  RECT 1376.460 0.000 1377.580 1.120 ;
  LAYER ME1 ;
  RECT 1376.460 0.000 1377.580 1.120 ;
 END
END DO91
PIN DI91
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1368.400 0.000 1369.520 1.120 ;
  LAYER ME3 ;
  RECT 1368.400 0.000 1369.520 1.120 ;
  LAYER ME2 ;
  RECT 1368.400 0.000 1369.520 1.120 ;
  LAYER ME1 ;
  RECT 1368.400 0.000 1369.520 1.120 ;
 END
END DI91
PIN DO90
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1363.440 0.000 1364.560 1.120 ;
  LAYER ME3 ;
  RECT 1363.440 0.000 1364.560 1.120 ;
  LAYER ME2 ;
  RECT 1363.440 0.000 1364.560 1.120 ;
  LAYER ME1 ;
  RECT 1363.440 0.000 1364.560 1.120 ;
 END
END DO90
PIN DI90
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1354.760 0.000 1355.880 1.120 ;
  LAYER ME3 ;
  RECT 1354.760 0.000 1355.880 1.120 ;
  LAYER ME2 ;
  RECT 1354.760 0.000 1355.880 1.120 ;
  LAYER ME1 ;
  RECT 1354.760 0.000 1355.880 1.120 ;
 END
END DI90
PIN DO89
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1346.700 0.000 1347.820 1.120 ;
  LAYER ME3 ;
  RECT 1346.700 0.000 1347.820 1.120 ;
  LAYER ME2 ;
  RECT 1346.700 0.000 1347.820 1.120 ;
  LAYER ME1 ;
  RECT 1346.700 0.000 1347.820 1.120 ;
 END
END DO89
PIN DI89
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1338.020 0.000 1339.140 1.120 ;
  LAYER ME3 ;
  RECT 1338.020 0.000 1339.140 1.120 ;
  LAYER ME2 ;
  RECT 1338.020 0.000 1339.140 1.120 ;
  LAYER ME1 ;
  RECT 1338.020 0.000 1339.140 1.120 ;
 END
END DI89
PIN DO88
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1333.060 0.000 1334.180 1.120 ;
  LAYER ME3 ;
  RECT 1333.060 0.000 1334.180 1.120 ;
  LAYER ME2 ;
  RECT 1333.060 0.000 1334.180 1.120 ;
  LAYER ME1 ;
  RECT 1333.060 0.000 1334.180 1.120 ;
 END
END DO88
PIN DI88
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1325.000 0.000 1326.120 1.120 ;
  LAYER ME3 ;
  RECT 1325.000 0.000 1326.120 1.120 ;
  LAYER ME2 ;
  RECT 1325.000 0.000 1326.120 1.120 ;
  LAYER ME1 ;
  RECT 1325.000 0.000 1326.120 1.120 ;
 END
END DI88
PIN DO87
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1320.040 0.000 1321.160 1.120 ;
  LAYER ME3 ;
  RECT 1320.040 0.000 1321.160 1.120 ;
  LAYER ME2 ;
  RECT 1320.040 0.000 1321.160 1.120 ;
  LAYER ME1 ;
  RECT 1320.040 0.000 1321.160 1.120 ;
 END
END DO87
PIN DI87
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1311.980 0.000 1313.100 1.120 ;
  LAYER ME3 ;
  RECT 1311.980 0.000 1313.100 1.120 ;
  LAYER ME2 ;
  RECT 1311.980 0.000 1313.100 1.120 ;
  LAYER ME1 ;
  RECT 1311.980 0.000 1313.100 1.120 ;
 END
END DI87
PIN DO86
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1307.020 0.000 1308.140 1.120 ;
  LAYER ME3 ;
  RECT 1307.020 0.000 1308.140 1.120 ;
  LAYER ME2 ;
  RECT 1307.020 0.000 1308.140 1.120 ;
  LAYER ME1 ;
  RECT 1307.020 0.000 1308.140 1.120 ;
 END
END DO86
PIN DI86
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1298.340 0.000 1299.460 1.120 ;
  LAYER ME3 ;
  RECT 1298.340 0.000 1299.460 1.120 ;
  LAYER ME2 ;
  RECT 1298.340 0.000 1299.460 1.120 ;
  LAYER ME1 ;
  RECT 1298.340 0.000 1299.460 1.120 ;
 END
END DI86
PIN DO85
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1290.280 0.000 1291.400 1.120 ;
  LAYER ME3 ;
  RECT 1290.280 0.000 1291.400 1.120 ;
  LAYER ME2 ;
  RECT 1290.280 0.000 1291.400 1.120 ;
  LAYER ME1 ;
  RECT 1290.280 0.000 1291.400 1.120 ;
 END
END DO85
PIN DI85
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1281.600 0.000 1282.720 1.120 ;
  LAYER ME3 ;
  RECT 1281.600 0.000 1282.720 1.120 ;
  LAYER ME2 ;
  RECT 1281.600 0.000 1282.720 1.120 ;
  LAYER ME1 ;
  RECT 1281.600 0.000 1282.720 1.120 ;
 END
END DI85
PIN DO84
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1276.640 0.000 1277.760 1.120 ;
  LAYER ME3 ;
  RECT 1276.640 0.000 1277.760 1.120 ;
  LAYER ME2 ;
  RECT 1276.640 0.000 1277.760 1.120 ;
  LAYER ME1 ;
  RECT 1276.640 0.000 1277.760 1.120 ;
 END
END DO84
PIN DI84
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1268.580 0.000 1269.700 1.120 ;
  LAYER ME3 ;
  RECT 1268.580 0.000 1269.700 1.120 ;
  LAYER ME2 ;
  RECT 1268.580 0.000 1269.700 1.120 ;
  LAYER ME1 ;
  RECT 1268.580 0.000 1269.700 1.120 ;
 END
END DI84
PIN DO83
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1263.620 0.000 1264.740 1.120 ;
  LAYER ME3 ;
  RECT 1263.620 0.000 1264.740 1.120 ;
  LAYER ME2 ;
  RECT 1263.620 0.000 1264.740 1.120 ;
  LAYER ME1 ;
  RECT 1263.620 0.000 1264.740 1.120 ;
 END
END DO83
PIN DI83
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1254.940 0.000 1256.060 1.120 ;
  LAYER ME3 ;
  RECT 1254.940 0.000 1256.060 1.120 ;
  LAYER ME2 ;
  RECT 1254.940 0.000 1256.060 1.120 ;
  LAYER ME1 ;
  RECT 1254.940 0.000 1256.060 1.120 ;
 END
END DI83
PIN DO82
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1249.980 0.000 1251.100 1.120 ;
  LAYER ME3 ;
  RECT 1249.980 0.000 1251.100 1.120 ;
  LAYER ME2 ;
  RECT 1249.980 0.000 1251.100 1.120 ;
  LAYER ME1 ;
  RECT 1249.980 0.000 1251.100 1.120 ;
 END
END DO82
PIN DI82
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1241.920 0.000 1243.040 1.120 ;
  LAYER ME3 ;
  RECT 1241.920 0.000 1243.040 1.120 ;
  LAYER ME2 ;
  RECT 1241.920 0.000 1243.040 1.120 ;
  LAYER ME1 ;
  RECT 1241.920 0.000 1243.040 1.120 ;
 END
END DI82
PIN DO81
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1233.860 0.000 1234.980 1.120 ;
  LAYER ME3 ;
  RECT 1233.860 0.000 1234.980 1.120 ;
  LAYER ME2 ;
  RECT 1233.860 0.000 1234.980 1.120 ;
  LAYER ME1 ;
  RECT 1233.860 0.000 1234.980 1.120 ;
 END
END DO81
PIN DI81
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1225.180 0.000 1226.300 1.120 ;
  LAYER ME3 ;
  RECT 1225.180 0.000 1226.300 1.120 ;
  LAYER ME2 ;
  RECT 1225.180 0.000 1226.300 1.120 ;
  LAYER ME1 ;
  RECT 1225.180 0.000 1226.300 1.120 ;
 END
END DI81
PIN DO80
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1220.220 0.000 1221.340 1.120 ;
  LAYER ME3 ;
  RECT 1220.220 0.000 1221.340 1.120 ;
  LAYER ME2 ;
  RECT 1220.220 0.000 1221.340 1.120 ;
  LAYER ME1 ;
  RECT 1220.220 0.000 1221.340 1.120 ;
 END
END DO80
PIN DI80
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1212.160 0.000 1213.280 1.120 ;
  LAYER ME3 ;
  RECT 1212.160 0.000 1213.280 1.120 ;
  LAYER ME2 ;
  RECT 1212.160 0.000 1213.280 1.120 ;
  LAYER ME1 ;
  RECT 1212.160 0.000 1213.280 1.120 ;
 END
END DI80
PIN DO79
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1207.200 0.000 1208.320 1.120 ;
  LAYER ME3 ;
  RECT 1207.200 0.000 1208.320 1.120 ;
  LAYER ME2 ;
  RECT 1207.200 0.000 1208.320 1.120 ;
  LAYER ME1 ;
  RECT 1207.200 0.000 1208.320 1.120 ;
 END
END DO79
PIN DI79
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1198.520 0.000 1199.640 1.120 ;
  LAYER ME3 ;
  RECT 1198.520 0.000 1199.640 1.120 ;
  LAYER ME2 ;
  RECT 1198.520 0.000 1199.640 1.120 ;
  LAYER ME1 ;
  RECT 1198.520 0.000 1199.640 1.120 ;
 END
END DI79
PIN DO78
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1193.560 0.000 1194.680 1.120 ;
  LAYER ME3 ;
  RECT 1193.560 0.000 1194.680 1.120 ;
  LAYER ME2 ;
  RECT 1193.560 0.000 1194.680 1.120 ;
  LAYER ME1 ;
  RECT 1193.560 0.000 1194.680 1.120 ;
 END
END DO78
PIN DI78
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1185.500 0.000 1186.620 1.120 ;
  LAYER ME3 ;
  RECT 1185.500 0.000 1186.620 1.120 ;
  LAYER ME2 ;
  RECT 1185.500 0.000 1186.620 1.120 ;
  LAYER ME1 ;
  RECT 1185.500 0.000 1186.620 1.120 ;
 END
END DI78
PIN DO77
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1176.820 0.000 1177.940 1.120 ;
  LAYER ME3 ;
  RECT 1176.820 0.000 1177.940 1.120 ;
  LAYER ME2 ;
  RECT 1176.820 0.000 1177.940 1.120 ;
  LAYER ME1 ;
  RECT 1176.820 0.000 1177.940 1.120 ;
 END
END DO77
PIN DI77
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER ME3 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER ME2 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER ME1 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
 END
END DI77
PIN DO76
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1163.800 0.000 1164.920 1.120 ;
  LAYER ME3 ;
  RECT 1163.800 0.000 1164.920 1.120 ;
  LAYER ME2 ;
  RECT 1163.800 0.000 1164.920 1.120 ;
  LAYER ME1 ;
  RECT 1163.800 0.000 1164.920 1.120 ;
 END
END DO76
PIN DI76
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER ME3 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER ME2 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER ME1 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
 END
END DI76
PIN DO75
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1150.780 0.000 1151.900 1.120 ;
  LAYER ME3 ;
  RECT 1150.780 0.000 1151.900 1.120 ;
  LAYER ME2 ;
  RECT 1150.780 0.000 1151.900 1.120 ;
  LAYER ME1 ;
  RECT 1150.780 0.000 1151.900 1.120 ;
 END
END DO75
PIN DI75
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1142.100 0.000 1143.220 1.120 ;
  LAYER ME3 ;
  RECT 1142.100 0.000 1143.220 1.120 ;
  LAYER ME2 ;
  RECT 1142.100 0.000 1143.220 1.120 ;
  LAYER ME1 ;
  RECT 1142.100 0.000 1143.220 1.120 ;
 END
END DI75
PIN DO74
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1137.140 0.000 1138.260 1.120 ;
  LAYER ME3 ;
  RECT 1137.140 0.000 1138.260 1.120 ;
  LAYER ME2 ;
  RECT 1137.140 0.000 1138.260 1.120 ;
  LAYER ME1 ;
  RECT 1137.140 0.000 1138.260 1.120 ;
 END
END DO74
PIN DI74
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1129.080 0.000 1130.200 1.120 ;
  LAYER ME3 ;
  RECT 1129.080 0.000 1130.200 1.120 ;
  LAYER ME2 ;
  RECT 1129.080 0.000 1130.200 1.120 ;
  LAYER ME1 ;
  RECT 1129.080 0.000 1130.200 1.120 ;
 END
END DI74
PIN DO73
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1120.400 0.000 1121.520 1.120 ;
  LAYER ME3 ;
  RECT 1120.400 0.000 1121.520 1.120 ;
  LAYER ME2 ;
  RECT 1120.400 0.000 1121.520 1.120 ;
  LAYER ME1 ;
  RECT 1120.400 0.000 1121.520 1.120 ;
 END
END DO73
PIN DI73
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1112.340 0.000 1113.460 1.120 ;
  LAYER ME3 ;
  RECT 1112.340 0.000 1113.460 1.120 ;
  LAYER ME2 ;
  RECT 1112.340 0.000 1113.460 1.120 ;
  LAYER ME1 ;
  RECT 1112.340 0.000 1113.460 1.120 ;
 END
END DI73
PIN DO72
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1107.380 0.000 1108.500 1.120 ;
  LAYER ME3 ;
  RECT 1107.380 0.000 1108.500 1.120 ;
  LAYER ME2 ;
  RECT 1107.380 0.000 1108.500 1.120 ;
  LAYER ME1 ;
  RECT 1107.380 0.000 1108.500 1.120 ;
 END
END DO72
PIN DI72
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1098.700 0.000 1099.820 1.120 ;
  LAYER ME3 ;
  RECT 1098.700 0.000 1099.820 1.120 ;
  LAYER ME2 ;
  RECT 1098.700 0.000 1099.820 1.120 ;
  LAYER ME1 ;
  RECT 1098.700 0.000 1099.820 1.120 ;
 END
END DI72
PIN DO71
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1093.740 0.000 1094.860 1.120 ;
  LAYER ME3 ;
  RECT 1093.740 0.000 1094.860 1.120 ;
  LAYER ME2 ;
  RECT 1093.740 0.000 1094.860 1.120 ;
  LAYER ME1 ;
  RECT 1093.740 0.000 1094.860 1.120 ;
 END
END DO71
PIN DI71
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1085.680 0.000 1086.800 1.120 ;
  LAYER ME3 ;
  RECT 1085.680 0.000 1086.800 1.120 ;
  LAYER ME2 ;
  RECT 1085.680 0.000 1086.800 1.120 ;
  LAYER ME1 ;
  RECT 1085.680 0.000 1086.800 1.120 ;
 END
END DI71
PIN DO70
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1080.720 0.000 1081.840 1.120 ;
  LAYER ME3 ;
  RECT 1080.720 0.000 1081.840 1.120 ;
  LAYER ME2 ;
  RECT 1080.720 0.000 1081.840 1.120 ;
  LAYER ME1 ;
  RECT 1080.720 0.000 1081.840 1.120 ;
 END
END DO70
PIN DI70
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1072.040 0.000 1073.160 1.120 ;
  LAYER ME3 ;
  RECT 1072.040 0.000 1073.160 1.120 ;
  LAYER ME2 ;
  RECT 1072.040 0.000 1073.160 1.120 ;
  LAYER ME1 ;
  RECT 1072.040 0.000 1073.160 1.120 ;
 END
END DI70
PIN DO69
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1063.980 0.000 1065.100 1.120 ;
  LAYER ME3 ;
  RECT 1063.980 0.000 1065.100 1.120 ;
  LAYER ME2 ;
  RECT 1063.980 0.000 1065.100 1.120 ;
  LAYER ME1 ;
  RECT 1063.980 0.000 1065.100 1.120 ;
 END
END DO69
PIN DI69
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1055.920 0.000 1057.040 1.120 ;
  LAYER ME3 ;
  RECT 1055.920 0.000 1057.040 1.120 ;
  LAYER ME2 ;
  RECT 1055.920 0.000 1057.040 1.120 ;
  LAYER ME1 ;
  RECT 1055.920 0.000 1057.040 1.120 ;
 END
END DI69
PIN DO68
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1050.960 0.000 1052.080 1.120 ;
  LAYER ME3 ;
  RECT 1050.960 0.000 1052.080 1.120 ;
  LAYER ME2 ;
  RECT 1050.960 0.000 1052.080 1.120 ;
  LAYER ME1 ;
  RECT 1050.960 0.000 1052.080 1.120 ;
 END
END DO68
PIN DI68
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1042.280 0.000 1043.400 1.120 ;
  LAYER ME3 ;
  RECT 1042.280 0.000 1043.400 1.120 ;
  LAYER ME2 ;
  RECT 1042.280 0.000 1043.400 1.120 ;
  LAYER ME1 ;
  RECT 1042.280 0.000 1043.400 1.120 ;
 END
END DI68
PIN DO67
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1037.320 0.000 1038.440 1.120 ;
  LAYER ME3 ;
  RECT 1037.320 0.000 1038.440 1.120 ;
  LAYER ME2 ;
  RECT 1037.320 0.000 1038.440 1.120 ;
  LAYER ME1 ;
  RECT 1037.320 0.000 1038.440 1.120 ;
 END
END DO67
PIN DI67
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1029.260 0.000 1030.380 1.120 ;
  LAYER ME3 ;
  RECT 1029.260 0.000 1030.380 1.120 ;
  LAYER ME2 ;
  RECT 1029.260 0.000 1030.380 1.120 ;
  LAYER ME1 ;
  RECT 1029.260 0.000 1030.380 1.120 ;
 END
END DI67
PIN DO66
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1024.300 0.000 1025.420 1.120 ;
  LAYER ME3 ;
  RECT 1024.300 0.000 1025.420 1.120 ;
  LAYER ME2 ;
  RECT 1024.300 0.000 1025.420 1.120 ;
  LAYER ME1 ;
  RECT 1024.300 0.000 1025.420 1.120 ;
 END
END DO66
PIN DI66
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 1015.620 0.000 1016.740 1.120 ;
  LAYER ME3 ;
  RECT 1015.620 0.000 1016.740 1.120 ;
  LAYER ME2 ;
  RECT 1015.620 0.000 1016.740 1.120 ;
  LAYER ME1 ;
  RECT 1015.620 0.000 1016.740 1.120 ;
 END
END DI66
PIN DO65
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER ME3 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER ME2 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER ME1 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
 END
END DO65
PIN DI65
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 998.880 0.000 1000.000 1.120 ;
  LAYER ME3 ;
  RECT 998.880 0.000 1000.000 1.120 ;
  LAYER ME2 ;
  RECT 998.880 0.000 1000.000 1.120 ;
  LAYER ME1 ;
  RECT 998.880 0.000 1000.000 1.120 ;
 END
END DI65
PIN DO64
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER ME3 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER ME2 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER ME1 ;
  RECT 994.540 0.000 995.660 1.120 ;
 END
END DO64
PIN DI64
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 985.860 0.000 986.980 1.120 ;
  LAYER ME3 ;
  RECT 985.860 0.000 986.980 1.120 ;
  LAYER ME2 ;
  RECT 985.860 0.000 986.980 1.120 ;
  LAYER ME1 ;
  RECT 985.860 0.000 986.980 1.120 ;
 END
END DI64
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER ME3 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER ME2 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER ME1 ;
  RECT 980.280 0.000 981.400 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER ME3 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER ME2 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER ME1 ;
  RECT 978.420 0.000 979.540 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 973.460 0.000 974.580 1.120 ;
  LAYER ME3 ;
  RECT 973.460 0.000 974.580 1.120 ;
  LAYER ME2 ;
  RECT 973.460 0.000 974.580 1.120 ;
  LAYER ME1 ;
  RECT 973.460 0.000 974.580 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 971.600 0.000 972.720 1.120 ;
  LAYER ME3 ;
  RECT 971.600 0.000 972.720 1.120 ;
  LAYER ME2 ;
  RECT 971.600 0.000 972.720 1.120 ;
  LAYER ME1 ;
  RECT 971.600 0.000 972.720 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER ME3 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER ME2 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER ME1 ;
  RECT 949.900 0.000 951.020 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 946.800 0.000 947.920 1.120 ;
  LAYER ME3 ;
  RECT 946.800 0.000 947.920 1.120 ;
  LAYER ME2 ;
  RECT 946.800 0.000 947.920 1.120 ;
  LAYER ME1 ;
  RECT 946.800 0.000 947.920 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 944.940 0.000 946.060 1.120 ;
  LAYER ME3 ;
  RECT 944.940 0.000 946.060 1.120 ;
  LAYER ME2 ;
  RECT 944.940 0.000 946.060 1.120 ;
  LAYER ME1 ;
  RECT 944.940 0.000 946.060 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER ME3 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER ME2 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER ME1 ;
  RECT 940.600 0.000 941.720 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER ME3 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER ME2 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER ME1 ;
  RECT 933.160 0.000 934.280 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER ME3 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER ME2 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER ME1 ;
  RECT 930.060 0.000 931.180 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER ME3 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER ME2 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER ME1 ;
  RECT 922.000 0.000 923.120 1.120 ;
 END
END A6
PIN DO63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 910.840 0.000 911.960 1.120 ;
  LAYER ME3 ;
  RECT 910.840 0.000 911.960 1.120 ;
  LAYER ME2 ;
  RECT 910.840 0.000 911.960 1.120 ;
  LAYER ME1 ;
  RECT 910.840 0.000 911.960 1.120 ;
 END
END DO63
PIN DI63
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 902.780 0.000 903.900 1.120 ;
  LAYER ME3 ;
  RECT 902.780 0.000 903.900 1.120 ;
  LAYER ME2 ;
  RECT 902.780 0.000 903.900 1.120 ;
  LAYER ME1 ;
  RECT 902.780 0.000 903.900 1.120 ;
 END
END DI63
PIN DO62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 897.820 0.000 898.940 1.120 ;
  LAYER ME3 ;
  RECT 897.820 0.000 898.940 1.120 ;
  LAYER ME2 ;
  RECT 897.820 0.000 898.940 1.120 ;
  LAYER ME1 ;
  RECT 897.820 0.000 898.940 1.120 ;
 END
END DO62
PIN DI62
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 889.140 0.000 890.260 1.120 ;
  LAYER ME3 ;
  RECT 889.140 0.000 890.260 1.120 ;
  LAYER ME2 ;
  RECT 889.140 0.000 890.260 1.120 ;
  LAYER ME1 ;
  RECT 889.140 0.000 890.260 1.120 ;
 END
END DI62
PIN DO61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 881.080 0.000 882.200 1.120 ;
  LAYER ME3 ;
  RECT 881.080 0.000 882.200 1.120 ;
  LAYER ME2 ;
  RECT 881.080 0.000 882.200 1.120 ;
  LAYER ME1 ;
  RECT 881.080 0.000 882.200 1.120 ;
 END
END DO61
PIN DI61
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER ME3 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER ME2 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER ME1 ;
  RECT 873.020 0.000 874.140 1.120 ;
 END
END DI61
PIN DO60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 868.060 0.000 869.180 1.120 ;
  LAYER ME3 ;
  RECT 868.060 0.000 869.180 1.120 ;
  LAYER ME2 ;
  RECT 868.060 0.000 869.180 1.120 ;
  LAYER ME1 ;
  RECT 868.060 0.000 869.180 1.120 ;
 END
END DO60
PIN DI60
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME3 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME2 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME1 ;
  RECT 859.380 0.000 860.500 1.120 ;
 END
END DI60
PIN DO59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 854.420 0.000 855.540 1.120 ;
  LAYER ME3 ;
  RECT 854.420 0.000 855.540 1.120 ;
  LAYER ME2 ;
  RECT 854.420 0.000 855.540 1.120 ;
  LAYER ME1 ;
  RECT 854.420 0.000 855.540 1.120 ;
 END
END DO59
PIN DI59
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 846.360 0.000 847.480 1.120 ;
  LAYER ME3 ;
  RECT 846.360 0.000 847.480 1.120 ;
  LAYER ME2 ;
  RECT 846.360 0.000 847.480 1.120 ;
  LAYER ME1 ;
  RECT 846.360 0.000 847.480 1.120 ;
 END
END DI59
PIN DO58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 841.400 0.000 842.520 1.120 ;
  LAYER ME3 ;
  RECT 841.400 0.000 842.520 1.120 ;
  LAYER ME2 ;
  RECT 841.400 0.000 842.520 1.120 ;
  LAYER ME1 ;
  RECT 841.400 0.000 842.520 1.120 ;
 END
END DO58
PIN DI58
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER ME3 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER ME2 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER ME1 ;
  RECT 832.720 0.000 833.840 1.120 ;
 END
END DI58
PIN DO57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER ME3 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER ME2 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER ME1 ;
  RECT 824.660 0.000 825.780 1.120 ;
 END
END DO57
PIN DI57
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER ME3 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER ME2 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER ME1 ;
  RECT 815.980 0.000 817.100 1.120 ;
 END
END DI57
PIN DO56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER ME3 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER ME2 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER ME1 ;
  RECT 811.640 0.000 812.760 1.120 ;
 END
END DO56
PIN DI56
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER ME3 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER ME2 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER ME1 ;
  RECT 802.960 0.000 804.080 1.120 ;
 END
END DI56
PIN DO55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 798.000 0.000 799.120 1.120 ;
  LAYER ME3 ;
  RECT 798.000 0.000 799.120 1.120 ;
  LAYER ME2 ;
  RECT 798.000 0.000 799.120 1.120 ;
  LAYER ME1 ;
  RECT 798.000 0.000 799.120 1.120 ;
 END
END DO55
PIN DI55
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 789.940 0.000 791.060 1.120 ;
  LAYER ME3 ;
  RECT 789.940 0.000 791.060 1.120 ;
  LAYER ME2 ;
  RECT 789.940 0.000 791.060 1.120 ;
  LAYER ME1 ;
  RECT 789.940 0.000 791.060 1.120 ;
 END
END DI55
PIN DO54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 784.980 0.000 786.100 1.120 ;
  LAYER ME3 ;
  RECT 784.980 0.000 786.100 1.120 ;
  LAYER ME2 ;
  RECT 784.980 0.000 786.100 1.120 ;
  LAYER ME1 ;
  RECT 784.980 0.000 786.100 1.120 ;
 END
END DO54
PIN DI54
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 776.300 0.000 777.420 1.120 ;
  LAYER ME3 ;
  RECT 776.300 0.000 777.420 1.120 ;
  LAYER ME2 ;
  RECT 776.300 0.000 777.420 1.120 ;
  LAYER ME1 ;
  RECT 776.300 0.000 777.420 1.120 ;
 END
END DI54
PIN DO53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 768.240 0.000 769.360 1.120 ;
  LAYER ME3 ;
  RECT 768.240 0.000 769.360 1.120 ;
  LAYER ME2 ;
  RECT 768.240 0.000 769.360 1.120 ;
  LAYER ME1 ;
  RECT 768.240 0.000 769.360 1.120 ;
 END
END DO53
PIN DI53
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 759.560 0.000 760.680 1.120 ;
  LAYER ME3 ;
  RECT 759.560 0.000 760.680 1.120 ;
  LAYER ME2 ;
  RECT 759.560 0.000 760.680 1.120 ;
  LAYER ME1 ;
  RECT 759.560 0.000 760.680 1.120 ;
 END
END DI53
PIN DO52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 754.600 0.000 755.720 1.120 ;
  LAYER ME3 ;
  RECT 754.600 0.000 755.720 1.120 ;
  LAYER ME2 ;
  RECT 754.600 0.000 755.720 1.120 ;
  LAYER ME1 ;
  RECT 754.600 0.000 755.720 1.120 ;
 END
END DO52
PIN DI52
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 746.540 0.000 747.660 1.120 ;
  LAYER ME3 ;
  RECT 746.540 0.000 747.660 1.120 ;
  LAYER ME2 ;
  RECT 746.540 0.000 747.660 1.120 ;
  LAYER ME1 ;
  RECT 746.540 0.000 747.660 1.120 ;
 END
END DI52
PIN DO51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 741.580 0.000 742.700 1.120 ;
  LAYER ME3 ;
  RECT 741.580 0.000 742.700 1.120 ;
  LAYER ME2 ;
  RECT 741.580 0.000 742.700 1.120 ;
  LAYER ME1 ;
  RECT 741.580 0.000 742.700 1.120 ;
 END
END DO51
PIN DI51
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME3 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME2 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME1 ;
  RECT 732.900 0.000 734.020 1.120 ;
 END
END DI51
PIN DO50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 728.560 0.000 729.680 1.120 ;
  LAYER ME3 ;
  RECT 728.560 0.000 729.680 1.120 ;
  LAYER ME2 ;
  RECT 728.560 0.000 729.680 1.120 ;
  LAYER ME1 ;
  RECT 728.560 0.000 729.680 1.120 ;
 END
END DO50
PIN DI50
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 719.880 0.000 721.000 1.120 ;
  LAYER ME3 ;
  RECT 719.880 0.000 721.000 1.120 ;
  LAYER ME2 ;
  RECT 719.880 0.000 721.000 1.120 ;
  LAYER ME1 ;
  RECT 719.880 0.000 721.000 1.120 ;
 END
END DI50
PIN DO49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER ME3 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER ME2 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER ME1 ;
  RECT 711.820 0.000 712.940 1.120 ;
 END
END DO49
PIN DI49
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER ME3 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER ME2 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER ME1 ;
  RECT 703.140 0.000 704.260 1.120 ;
 END
END DI49
PIN DO48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER ME3 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER ME2 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER ME1 ;
  RECT 698.180 0.000 699.300 1.120 ;
 END
END DO48
PIN DI48
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER ME3 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER ME2 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER ME1 ;
  RECT 690.120 0.000 691.240 1.120 ;
 END
END DI48
PIN DO47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 685.160 0.000 686.280 1.120 ;
  LAYER ME3 ;
  RECT 685.160 0.000 686.280 1.120 ;
  LAYER ME2 ;
  RECT 685.160 0.000 686.280 1.120 ;
  LAYER ME1 ;
  RECT 685.160 0.000 686.280 1.120 ;
 END
END DO47
PIN DI47
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME3 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME2 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME1 ;
  RECT 676.480 0.000 677.600 1.120 ;
 END
END DI47
PIN DO46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER ME3 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER ME2 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER ME1 ;
  RECT 671.520 0.000 672.640 1.120 ;
 END
END DO46
PIN DI46
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 663.460 0.000 664.580 1.120 ;
  LAYER ME3 ;
  RECT 663.460 0.000 664.580 1.120 ;
  LAYER ME2 ;
  RECT 663.460 0.000 664.580 1.120 ;
  LAYER ME1 ;
  RECT 663.460 0.000 664.580 1.120 ;
 END
END DI46
PIN DO45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 654.780 0.000 655.900 1.120 ;
  LAYER ME3 ;
  RECT 654.780 0.000 655.900 1.120 ;
  LAYER ME2 ;
  RECT 654.780 0.000 655.900 1.120 ;
  LAYER ME1 ;
  RECT 654.780 0.000 655.900 1.120 ;
 END
END DO45
PIN DI45
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 646.720 0.000 647.840 1.120 ;
  LAYER ME3 ;
  RECT 646.720 0.000 647.840 1.120 ;
  LAYER ME2 ;
  RECT 646.720 0.000 647.840 1.120 ;
  LAYER ME1 ;
  RECT 646.720 0.000 647.840 1.120 ;
 END
END DI45
PIN DO44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME3 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME2 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME1 ;
  RECT 641.760 0.000 642.880 1.120 ;
 END
END DO44
PIN DI44
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME3 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME2 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME1 ;
  RECT 633.700 0.000 634.820 1.120 ;
 END
END DI44
PIN DO43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME3 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME2 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME1 ;
  RECT 628.740 0.000 629.860 1.120 ;
 END
END DO43
PIN DI43
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME3 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME2 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME1 ;
  RECT 620.060 0.000 621.180 1.120 ;
 END
END DI43
PIN DO42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 615.100 0.000 616.220 1.120 ;
  LAYER ME3 ;
  RECT 615.100 0.000 616.220 1.120 ;
  LAYER ME2 ;
  RECT 615.100 0.000 616.220 1.120 ;
  LAYER ME1 ;
  RECT 615.100 0.000 616.220 1.120 ;
 END
END DO42
PIN DI42
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 607.040 0.000 608.160 1.120 ;
  LAYER ME3 ;
  RECT 607.040 0.000 608.160 1.120 ;
  LAYER ME2 ;
  RECT 607.040 0.000 608.160 1.120 ;
  LAYER ME1 ;
  RECT 607.040 0.000 608.160 1.120 ;
 END
END DI42
PIN DO41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME3 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME2 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME1 ;
  RECT 598.360 0.000 599.480 1.120 ;
 END
END DO41
PIN DI41
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME3 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME2 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME1 ;
  RECT 590.300 0.000 591.420 1.120 ;
 END
END DI41
PIN DO40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME3 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME2 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME1 ;
  RECT 585.340 0.000 586.460 1.120 ;
 END
END DO40
PIN DI40
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME3 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME2 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME1 ;
  RECT 576.660 0.000 577.780 1.120 ;
 END
END DI40
PIN DO39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 571.700 0.000 572.820 1.120 ;
  LAYER ME3 ;
  RECT 571.700 0.000 572.820 1.120 ;
  LAYER ME2 ;
  RECT 571.700 0.000 572.820 1.120 ;
  LAYER ME1 ;
  RECT 571.700 0.000 572.820 1.120 ;
 END
END DO39
PIN DI39
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME3 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME2 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME1 ;
  RECT 563.640 0.000 564.760 1.120 ;
 END
END DI39
PIN DO38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 558.680 0.000 559.800 1.120 ;
  LAYER ME3 ;
  RECT 558.680 0.000 559.800 1.120 ;
  LAYER ME2 ;
  RECT 558.680 0.000 559.800 1.120 ;
  LAYER ME1 ;
  RECT 558.680 0.000 559.800 1.120 ;
 END
END DO38
PIN DI38
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER ME3 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER ME2 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER ME1 ;
  RECT 550.620 0.000 551.740 1.120 ;
 END
END DI38
PIN DO37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME3 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME2 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME1 ;
  RECT 541.940 0.000 543.060 1.120 ;
 END
END DO37
PIN DI37
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME3 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME2 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME1 ;
  RECT 533.880 0.000 535.000 1.120 ;
 END
END DI37
PIN DO36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME3 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME2 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME1 ;
  RECT 528.920 0.000 530.040 1.120 ;
 END
END DO36
PIN DI36
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME3 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME2 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME1 ;
  RECT 520.240 0.000 521.360 1.120 ;
 END
END DI36
PIN DO35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME3 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME2 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME1 ;
  RECT 515.280 0.000 516.400 1.120 ;
 END
END DO35
PIN DI35
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME3 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME2 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME1 ;
  RECT 507.220 0.000 508.340 1.120 ;
 END
END DI35
PIN DO34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 502.260 0.000 503.380 1.120 ;
  LAYER ME3 ;
  RECT 502.260 0.000 503.380 1.120 ;
  LAYER ME2 ;
  RECT 502.260 0.000 503.380 1.120 ;
  LAYER ME1 ;
  RECT 502.260 0.000 503.380 1.120 ;
 END
END DO34
PIN DI34
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 493.580 0.000 494.700 1.120 ;
  LAYER ME3 ;
  RECT 493.580 0.000 494.700 1.120 ;
  LAYER ME2 ;
  RECT 493.580 0.000 494.700 1.120 ;
  LAYER ME1 ;
  RECT 493.580 0.000 494.700 1.120 ;
 END
END DI34
PIN DO33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME3 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME2 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME1 ;
  RECT 485.520 0.000 486.640 1.120 ;
 END
END DO33
PIN DI33
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER ME3 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER ME2 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER ME1 ;
  RECT 476.840 0.000 477.960 1.120 ;
 END
END DI33
PIN DO32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME3 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME2 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME1 ;
  RECT 472.500 0.000 473.620 1.120 ;
 END
END DO32
PIN DI32
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME3 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME2 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME1 ;
  RECT 463.820 0.000 464.940 1.120 ;
 END
END DI32
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME3 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME2 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME1 ;
  RECT 458.860 0.000 459.980 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME3 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME2 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME1 ;
  RECT 450.800 0.000 451.920 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER ME3 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER ME2 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER ME1 ;
  RECT 445.840 0.000 446.960 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER ME3 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER ME2 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER ME1 ;
  RECT 437.160 0.000 438.280 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME3 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME2 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME1 ;
  RECT 420.420 0.000 421.540 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME3 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME2 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME1 ;
  RECT 415.460 0.000 416.580 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME3 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME2 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME1 ;
  RECT 407.400 0.000 408.520 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER ME3 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER ME2 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER ME1 ;
  RECT 393.760 0.000 394.880 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER ME3 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER ME2 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER ME1 ;
  RECT 389.420 0.000 390.540 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER ME3 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER ME2 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER ME1 ;
  RECT 380.740 0.000 381.860 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME3 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME2 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME1 ;
  RECT 372.680 0.000 373.800 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME3 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME2 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME1 ;
  RECT 364.000 0.000 365.120 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME3 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME2 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME1 ;
  RECT 350.980 0.000 352.100 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME3 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME2 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME1 ;
  RECT 346.020 0.000 347.140 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME3 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME2 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME1 ;
  RECT 337.340 0.000 338.460 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME3 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME2 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME1 ;
  RECT 332.380 0.000 333.500 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER ME3 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER ME2 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER ME1 ;
  RECT 324.320 0.000 325.440 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME3 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME2 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME1 ;
  RECT 316.260 0.000 317.380 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME3 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME2 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME1 ;
  RECT 307.580 0.000 308.700 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME3 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME2 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME1 ;
  RECT 302.620 0.000 303.740 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME3 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME2 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME1 ;
  RECT 294.560 0.000 295.680 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME3 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME2 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME1 ;
  RECT 280.920 0.000 282.040 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME3 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME2 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME1 ;
  RECT 275.960 0.000 277.080 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI16
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 1899.060 176.400 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 1899.060 176.400 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 1899.060 176.400 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 1899.060 176.400 ;
  LAYER VI1 ;
  RECT 0.000 0.140 1899.060 176.400 ;
  LAYER VI2 ;
  RECT 0.000 0.140 1899.060 176.400 ;
  LAYER VI3 ;
  RECT 0.000 0.140 1899.060 176.400 ;
END
END MID_SRAM.v
END LIBRARY



