# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SUMA180_256X16
#       Words            : 256
#       Bits             : 16
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2025/06/05 11:31:30
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SUMA180_256X16
CLASS BLOCK ;
FOREIGN SUMA180_256X16 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 316.200 BY 215.600 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 315.080 204.180 316.200 207.420 ;
  LAYER ME3 ;
  RECT 315.080 204.180 316.200 207.420 ;
  LAYER ME2 ;
  RECT 315.080 204.180 316.200 207.420 ;
  LAYER ME1 ;
  RECT 315.080 204.180 316.200 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 196.340 316.200 199.580 ;
  LAYER ME3 ;
  RECT 315.080 196.340 316.200 199.580 ;
  LAYER ME2 ;
  RECT 315.080 196.340 316.200 199.580 ;
  LAYER ME1 ;
  RECT 315.080 196.340 316.200 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 188.500 316.200 191.740 ;
  LAYER ME3 ;
  RECT 315.080 188.500 316.200 191.740 ;
  LAYER ME2 ;
  RECT 315.080 188.500 316.200 191.740 ;
  LAYER ME1 ;
  RECT 315.080 188.500 316.200 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 180.660 316.200 183.900 ;
  LAYER ME3 ;
  RECT 315.080 180.660 316.200 183.900 ;
  LAYER ME2 ;
  RECT 315.080 180.660 316.200 183.900 ;
  LAYER ME1 ;
  RECT 315.080 180.660 316.200 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 172.820 316.200 176.060 ;
  LAYER ME3 ;
  RECT 315.080 172.820 316.200 176.060 ;
  LAYER ME2 ;
  RECT 315.080 172.820 316.200 176.060 ;
  LAYER ME1 ;
  RECT 315.080 172.820 316.200 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 164.980 316.200 168.220 ;
  LAYER ME3 ;
  RECT 315.080 164.980 316.200 168.220 ;
  LAYER ME2 ;
  RECT 315.080 164.980 316.200 168.220 ;
  LAYER ME1 ;
  RECT 315.080 164.980 316.200 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 125.780 316.200 129.020 ;
  LAYER ME3 ;
  RECT 315.080 125.780 316.200 129.020 ;
  LAYER ME2 ;
  RECT 315.080 125.780 316.200 129.020 ;
  LAYER ME1 ;
  RECT 315.080 125.780 316.200 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 117.940 316.200 121.180 ;
  LAYER ME3 ;
  RECT 315.080 117.940 316.200 121.180 ;
  LAYER ME2 ;
  RECT 315.080 117.940 316.200 121.180 ;
  LAYER ME1 ;
  RECT 315.080 117.940 316.200 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 110.100 316.200 113.340 ;
  LAYER ME3 ;
  RECT 315.080 110.100 316.200 113.340 ;
  LAYER ME2 ;
  RECT 315.080 110.100 316.200 113.340 ;
  LAYER ME1 ;
  RECT 315.080 110.100 316.200 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 102.260 316.200 105.500 ;
  LAYER ME3 ;
  RECT 315.080 102.260 316.200 105.500 ;
  LAYER ME2 ;
  RECT 315.080 102.260 316.200 105.500 ;
  LAYER ME1 ;
  RECT 315.080 102.260 316.200 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 94.420 316.200 97.660 ;
  LAYER ME3 ;
  RECT 315.080 94.420 316.200 97.660 ;
  LAYER ME2 ;
  RECT 315.080 94.420 316.200 97.660 ;
  LAYER ME1 ;
  RECT 315.080 94.420 316.200 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 86.580 316.200 89.820 ;
  LAYER ME3 ;
  RECT 315.080 86.580 316.200 89.820 ;
  LAYER ME2 ;
  RECT 315.080 86.580 316.200 89.820 ;
  LAYER ME1 ;
  RECT 315.080 86.580 316.200 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 47.380 316.200 50.620 ;
  LAYER ME3 ;
  RECT 315.080 47.380 316.200 50.620 ;
  LAYER ME2 ;
  RECT 315.080 47.380 316.200 50.620 ;
  LAYER ME1 ;
  RECT 315.080 47.380 316.200 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 39.540 316.200 42.780 ;
  LAYER ME3 ;
  RECT 315.080 39.540 316.200 42.780 ;
  LAYER ME2 ;
  RECT 315.080 39.540 316.200 42.780 ;
  LAYER ME1 ;
  RECT 315.080 39.540 316.200 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 31.700 316.200 34.940 ;
  LAYER ME3 ;
  RECT 315.080 31.700 316.200 34.940 ;
  LAYER ME2 ;
  RECT 315.080 31.700 316.200 34.940 ;
  LAYER ME1 ;
  RECT 315.080 31.700 316.200 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 23.860 316.200 27.100 ;
  LAYER ME3 ;
  RECT 315.080 23.860 316.200 27.100 ;
  LAYER ME2 ;
  RECT 315.080 23.860 316.200 27.100 ;
  LAYER ME1 ;
  RECT 315.080 23.860 316.200 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 16.020 316.200 19.260 ;
  LAYER ME3 ;
  RECT 315.080 16.020 316.200 19.260 ;
  LAYER ME2 ;
  RECT 315.080 16.020 316.200 19.260 ;
  LAYER ME1 ;
  RECT 315.080 16.020 316.200 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 8.180 316.200 11.420 ;
  LAYER ME3 ;
  RECT 315.080 8.180 316.200 11.420 ;
  LAYER ME2 ;
  RECT 315.080 8.180 316.200 11.420 ;
  LAYER ME1 ;
  RECT 315.080 8.180 316.200 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 214.480 306.500 215.600 ;
  LAYER ME3 ;
  RECT 302.960 214.480 306.500 215.600 ;
  LAYER ME2 ;
  RECT 302.960 214.480 306.500 215.600 ;
  LAYER ME1 ;
  RECT 302.960 214.480 306.500 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 214.480 297.820 215.600 ;
  LAYER ME3 ;
  RECT 294.280 214.480 297.820 215.600 ;
  LAYER ME2 ;
  RECT 294.280 214.480 297.820 215.600 ;
  LAYER ME1 ;
  RECT 294.280 214.480 297.820 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 214.480 289.140 215.600 ;
  LAYER ME3 ;
  RECT 285.600 214.480 289.140 215.600 ;
  LAYER ME2 ;
  RECT 285.600 214.480 289.140 215.600 ;
  LAYER ME1 ;
  RECT 285.600 214.480 289.140 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 214.480 280.460 215.600 ;
  LAYER ME3 ;
  RECT 276.920 214.480 280.460 215.600 ;
  LAYER ME2 ;
  RECT 276.920 214.480 280.460 215.600 ;
  LAYER ME1 ;
  RECT 276.920 214.480 280.460 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 214.480 271.780 215.600 ;
  LAYER ME3 ;
  RECT 268.240 214.480 271.780 215.600 ;
  LAYER ME2 ;
  RECT 268.240 214.480 271.780 215.600 ;
  LAYER ME1 ;
  RECT 268.240 214.480 271.780 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 214.480 228.380 215.600 ;
  LAYER ME3 ;
  RECT 224.840 214.480 228.380 215.600 ;
  LAYER ME2 ;
  RECT 224.840 214.480 228.380 215.600 ;
  LAYER ME1 ;
  RECT 224.840 214.480 228.380 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 214.480 219.700 215.600 ;
  LAYER ME3 ;
  RECT 216.160 214.480 219.700 215.600 ;
  LAYER ME2 ;
  RECT 216.160 214.480 219.700 215.600 ;
  LAYER ME1 ;
  RECT 216.160 214.480 219.700 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 214.480 211.020 215.600 ;
  LAYER ME3 ;
  RECT 207.480 214.480 211.020 215.600 ;
  LAYER ME2 ;
  RECT 207.480 214.480 211.020 215.600 ;
  LAYER ME1 ;
  RECT 207.480 214.480 211.020 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 214.480 202.340 215.600 ;
  LAYER ME3 ;
  RECT 198.800 214.480 202.340 215.600 ;
  LAYER ME2 ;
  RECT 198.800 214.480 202.340 215.600 ;
  LAYER ME1 ;
  RECT 198.800 214.480 202.340 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER ME3 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER ME2 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER ME1 ;
  RECT 190.120 214.480 193.660 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER ME3 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER ME2 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER ME1 ;
  RECT 181.440 214.480 184.980 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER ME3 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER ME2 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER ME1 ;
  RECT 138.040 214.480 141.580 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER ME3 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER ME2 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER ME1 ;
  RECT 129.360 214.480 132.900 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER ME3 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER ME2 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER ME1 ;
  RECT 120.680 214.480 124.220 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER ME3 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER ME2 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER ME1 ;
  RECT 112.000 214.480 115.540 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER ME3 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER ME2 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER ME1 ;
  RECT 103.320 214.480 106.860 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER ME3 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER ME2 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER ME1 ;
  RECT 94.640 214.480 98.180 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER ME3 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER ME2 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER ME1 ;
  RECT 51.240 214.480 54.780 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER ME3 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER ME2 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER ME1 ;
  RECT 42.560 214.480 46.100 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER ME3 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER ME2 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER ME1 ;
  RECT 33.880 214.480 37.420 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER ME3 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER ME2 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER ME1 ;
  RECT 25.200 214.480 28.740 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER ME3 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER ME2 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER ME1 ;
  RECT 16.520 214.480 20.060 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER ME3 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER ME2 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER ME1 ;
  RECT 7.840 214.480 11.380 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME3 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME2 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME1 ;
  RECT 296.760 0.000 300.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.060 0.000 278.600 1.120 ;
  LAYER ME3 ;
  RECT 275.060 0.000 278.600 1.120 ;
  LAYER ME2 ;
  RECT 275.060 0.000 278.600 1.120 ;
  LAYER ME1 ;
  RECT 275.060 0.000 278.600 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER ME3 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER ME2 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER ME1 ;
  RECT 226.700 0.000 230.240 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME3 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME2 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME1 ;
  RECT 121.920 0.000 125.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 315.080 200.260 316.200 203.500 ;
  LAYER ME3 ;
  RECT 315.080 200.260 316.200 203.500 ;
  LAYER ME2 ;
  RECT 315.080 200.260 316.200 203.500 ;
  LAYER ME1 ;
  RECT 315.080 200.260 316.200 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 192.420 316.200 195.660 ;
  LAYER ME3 ;
  RECT 315.080 192.420 316.200 195.660 ;
  LAYER ME2 ;
  RECT 315.080 192.420 316.200 195.660 ;
  LAYER ME1 ;
  RECT 315.080 192.420 316.200 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 184.580 316.200 187.820 ;
  LAYER ME3 ;
  RECT 315.080 184.580 316.200 187.820 ;
  LAYER ME2 ;
  RECT 315.080 184.580 316.200 187.820 ;
  LAYER ME1 ;
  RECT 315.080 184.580 316.200 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 176.740 316.200 179.980 ;
  LAYER ME3 ;
  RECT 315.080 176.740 316.200 179.980 ;
  LAYER ME2 ;
  RECT 315.080 176.740 316.200 179.980 ;
  LAYER ME1 ;
  RECT 315.080 176.740 316.200 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 168.900 316.200 172.140 ;
  LAYER ME3 ;
  RECT 315.080 168.900 316.200 172.140 ;
  LAYER ME2 ;
  RECT 315.080 168.900 316.200 172.140 ;
  LAYER ME1 ;
  RECT 315.080 168.900 316.200 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 129.700 316.200 132.940 ;
  LAYER ME3 ;
  RECT 315.080 129.700 316.200 132.940 ;
  LAYER ME2 ;
  RECT 315.080 129.700 316.200 132.940 ;
  LAYER ME1 ;
  RECT 315.080 129.700 316.200 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 121.860 316.200 125.100 ;
  LAYER ME3 ;
  RECT 315.080 121.860 316.200 125.100 ;
  LAYER ME2 ;
  RECT 315.080 121.860 316.200 125.100 ;
  LAYER ME1 ;
  RECT 315.080 121.860 316.200 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 114.020 316.200 117.260 ;
  LAYER ME3 ;
  RECT 315.080 114.020 316.200 117.260 ;
  LAYER ME2 ;
  RECT 315.080 114.020 316.200 117.260 ;
  LAYER ME1 ;
  RECT 315.080 114.020 316.200 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 106.180 316.200 109.420 ;
  LAYER ME3 ;
  RECT 315.080 106.180 316.200 109.420 ;
  LAYER ME2 ;
  RECT 315.080 106.180 316.200 109.420 ;
  LAYER ME1 ;
  RECT 315.080 106.180 316.200 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 98.340 316.200 101.580 ;
  LAYER ME3 ;
  RECT 315.080 98.340 316.200 101.580 ;
  LAYER ME2 ;
  RECT 315.080 98.340 316.200 101.580 ;
  LAYER ME1 ;
  RECT 315.080 98.340 316.200 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 90.500 316.200 93.740 ;
  LAYER ME3 ;
  RECT 315.080 90.500 316.200 93.740 ;
  LAYER ME2 ;
  RECT 315.080 90.500 316.200 93.740 ;
  LAYER ME1 ;
  RECT 315.080 90.500 316.200 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 51.300 316.200 54.540 ;
  LAYER ME3 ;
  RECT 315.080 51.300 316.200 54.540 ;
  LAYER ME2 ;
  RECT 315.080 51.300 316.200 54.540 ;
  LAYER ME1 ;
  RECT 315.080 51.300 316.200 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 43.460 316.200 46.700 ;
  LAYER ME3 ;
  RECT 315.080 43.460 316.200 46.700 ;
  LAYER ME2 ;
  RECT 315.080 43.460 316.200 46.700 ;
  LAYER ME1 ;
  RECT 315.080 43.460 316.200 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 35.620 316.200 38.860 ;
  LAYER ME3 ;
  RECT 315.080 35.620 316.200 38.860 ;
  LAYER ME2 ;
  RECT 315.080 35.620 316.200 38.860 ;
  LAYER ME1 ;
  RECT 315.080 35.620 316.200 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 27.780 316.200 31.020 ;
  LAYER ME3 ;
  RECT 315.080 27.780 316.200 31.020 ;
  LAYER ME2 ;
  RECT 315.080 27.780 316.200 31.020 ;
  LAYER ME1 ;
  RECT 315.080 27.780 316.200 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 19.940 316.200 23.180 ;
  LAYER ME3 ;
  RECT 315.080 19.940 316.200 23.180 ;
  LAYER ME2 ;
  RECT 315.080 19.940 316.200 23.180 ;
  LAYER ME1 ;
  RECT 315.080 19.940 316.200 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.080 12.100 316.200 15.340 ;
  LAYER ME3 ;
  RECT 315.080 12.100 316.200 15.340 ;
  LAYER ME2 ;
  RECT 315.080 12.100 316.200 15.340 ;
  LAYER ME1 ;
  RECT 315.080 12.100 316.200 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 214.480 302.160 215.600 ;
  LAYER ME3 ;
  RECT 298.620 214.480 302.160 215.600 ;
  LAYER ME2 ;
  RECT 298.620 214.480 302.160 215.600 ;
  LAYER ME1 ;
  RECT 298.620 214.480 302.160 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 214.480 293.480 215.600 ;
  LAYER ME3 ;
  RECT 289.940 214.480 293.480 215.600 ;
  LAYER ME2 ;
  RECT 289.940 214.480 293.480 215.600 ;
  LAYER ME1 ;
  RECT 289.940 214.480 293.480 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 214.480 284.800 215.600 ;
  LAYER ME3 ;
  RECT 281.260 214.480 284.800 215.600 ;
  LAYER ME2 ;
  RECT 281.260 214.480 284.800 215.600 ;
  LAYER ME1 ;
  RECT 281.260 214.480 284.800 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 214.480 276.120 215.600 ;
  LAYER ME3 ;
  RECT 272.580 214.480 276.120 215.600 ;
  LAYER ME2 ;
  RECT 272.580 214.480 276.120 215.600 ;
  LAYER ME1 ;
  RECT 272.580 214.480 276.120 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 214.480 232.720 215.600 ;
  LAYER ME3 ;
  RECT 229.180 214.480 232.720 215.600 ;
  LAYER ME2 ;
  RECT 229.180 214.480 232.720 215.600 ;
  LAYER ME1 ;
  RECT 229.180 214.480 232.720 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 214.480 224.040 215.600 ;
  LAYER ME3 ;
  RECT 220.500 214.480 224.040 215.600 ;
  LAYER ME2 ;
  RECT 220.500 214.480 224.040 215.600 ;
  LAYER ME1 ;
  RECT 220.500 214.480 224.040 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 214.480 215.360 215.600 ;
  LAYER ME3 ;
  RECT 211.820 214.480 215.360 215.600 ;
  LAYER ME2 ;
  RECT 211.820 214.480 215.360 215.600 ;
  LAYER ME1 ;
  RECT 211.820 214.480 215.360 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 214.480 206.680 215.600 ;
  LAYER ME3 ;
  RECT 203.140 214.480 206.680 215.600 ;
  LAYER ME2 ;
  RECT 203.140 214.480 206.680 215.600 ;
  LAYER ME1 ;
  RECT 203.140 214.480 206.680 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 214.480 198.000 215.600 ;
  LAYER ME3 ;
  RECT 194.460 214.480 198.000 215.600 ;
  LAYER ME2 ;
  RECT 194.460 214.480 198.000 215.600 ;
  LAYER ME1 ;
  RECT 194.460 214.480 198.000 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER ME3 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER ME2 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER ME1 ;
  RECT 185.780 214.480 189.320 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER ME3 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER ME2 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER ME1 ;
  RECT 142.380 214.480 145.920 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER ME3 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER ME2 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER ME1 ;
  RECT 133.700 214.480 137.240 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER ME3 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER ME2 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER ME1 ;
  RECT 125.020 214.480 128.560 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER ME3 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER ME2 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER ME1 ;
  RECT 116.340 214.480 119.880 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER ME3 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER ME2 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER ME1 ;
  RECT 107.660 214.480 111.200 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER ME3 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER ME2 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER ME1 ;
  RECT 98.980 214.480 102.520 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER ME3 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER ME2 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER ME1 ;
  RECT 55.580 214.480 59.120 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER ME3 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER ME2 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER ME1 ;
  RECT 46.900 214.480 50.440 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER ME3 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER ME2 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER ME1 ;
  RECT 38.220 214.480 41.760 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER ME3 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER ME2 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER ME1 ;
  RECT 29.540 214.480 33.080 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER ME3 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER ME2 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER ME1 ;
  RECT 20.860 214.480 24.400 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER ME3 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER ME2 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER ME1 ;
  RECT 12.180 214.480 15.720 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER ME3 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER ME2 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER ME1 ;
  RECT 304.820 0.000 308.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 266.380 0.000 269.920 1.120 ;
  LAYER ME3 ;
  RECT 266.380 0.000 269.920 1.120 ;
  LAYER ME2 ;
  RECT 266.380 0.000 269.920 1.120 ;
  LAYER ME1 ;
  RECT 266.380 0.000 269.920 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER ME3 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER ME2 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER ME1 ;
  RECT 133.080 0.000 136.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME3 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME2 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME1 ;
  RECT 302.620 0.000 303.740 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME3 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME2 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME1 ;
  RECT 294.560 0.000 295.680 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME3 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME2 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME1 ;
  RECT 280.920 0.000 282.040 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER ME3 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER ME2 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER ME1 ;
  RECT 272.860 0.000 273.980 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 264.180 0.000 265.300 1.120 ;
  LAYER ME3 ;
  RECT 264.180 0.000 265.300 1.120 ;
  LAYER ME2 ;
  RECT 264.180 0.000 265.300 1.120 ;
  LAYER ME1 ;
  RECT 264.180 0.000 265.300 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 216.440 0.000 217.560 1.120 ;
  LAYER ME3 ;
  RECT 216.440 0.000 217.560 1.120 ;
  LAYER ME2 ;
  RECT 216.440 0.000 217.560 1.120 ;
  LAYER ME1 ;
  RECT 216.440 0.000 217.560 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 207.760 0.000 208.880 1.120 ;
  LAYER ME3 ;
  RECT 207.760 0.000 208.880 1.120 ;
  LAYER ME2 ;
  RECT 207.760 0.000 208.880 1.120 ;
  LAYER ME1 ;
  RECT 207.760 0.000 208.880 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI8
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 189.160 0.000 190.280 1.120 ;
  LAYER ME3 ;
  RECT 189.160 0.000 190.280 1.120 ;
  LAYER ME2 ;
  RECT 189.160 0.000 190.280 1.120 ;
  LAYER ME1 ;
  RECT 189.160 0.000 190.280 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER ME3 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER ME2 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER ME1 ;
  RECT 182.340 0.000 183.460 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 180.480 0.000 181.600 1.120 ;
  LAYER ME3 ;
  RECT 180.480 0.000 181.600 1.120 ;
  LAYER ME2 ;
  RECT 180.480 0.000 181.600 1.120 ;
  LAYER ME1 ;
  RECT 180.480 0.000 181.600 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 158.780 0.000 159.900 1.120 ;
  LAYER ME3 ;
  RECT 158.780 0.000 159.900 1.120 ;
  LAYER ME2 ;
  RECT 158.780 0.000 159.900 1.120 ;
  LAYER ME1 ;
  RECT 158.780 0.000 159.900 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 155.680 0.000 156.800 1.120 ;
  LAYER ME3 ;
  RECT 155.680 0.000 156.800 1.120 ;
  LAYER ME2 ;
  RECT 155.680 0.000 156.800 1.120 ;
  LAYER ME1 ;
  RECT 155.680 0.000 156.800 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 153.200 0.000 154.320 1.120 ;
  LAYER ME3 ;
  RECT 153.200 0.000 154.320 1.120 ;
  LAYER ME2 ;
  RECT 153.200 0.000 154.320 1.120 ;
  LAYER ME1 ;
  RECT 153.200 0.000 154.320 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME3 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME2 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME1 ;
  RECT 148.860 0.000 149.980 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME3 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME2 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME1 ;
  RECT 141.420 0.000 142.540 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME3 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME2 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME1 ;
  RECT 138.320 0.000 139.440 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME3 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME2 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME1 ;
  RECT 130.880 0.000 132.000 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER ME3 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER ME2 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER ME1 ;
  RECT 127.780 0.000 128.900 1.120 ;
 END
END A7
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 316.200 215.600 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 316.200 215.600 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 316.200 215.600 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 316.200 215.600 ;
  LAYER VI1 ;
  RECT 0.000 0.140 316.200 215.600 ;
  LAYER VI2 ;
  RECT 0.000 0.140 316.200 215.600 ;
  LAYER VI3 ;
  RECT 0.000 0.140 316.200 215.600 ;
END
END SUMA180_256X16
END LIBRARY



