/RAID2/COURSE/iclab/iclabTA07/DemoEnv_2025/01_RTL/AFS.sv