../00_TESTBED/INF.sv