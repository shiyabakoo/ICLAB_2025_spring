//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab04 Exercise		: Two Head Attention
//   Author     		: Yu-Chi Lin (a6121461214.st12@nycu.edu.tw)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : ATTN.v
//   Module Name : ATTN
//   Release version : V1.0 (Release Date: 2025-3)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME      50.0
`define SEED_NUMBER     28825252
`define PATTERN_NUMBER 100

module PATTERN
`protected
2S.M8P<VH<^SS>9eAQV[D8a?>M]PbQ@49.aa#W0<?=53L5ZM9W9R&)LIa247OeD0
,GZEad?QdEHP]_N4W-cc<^\SdV:S0<\9MZG3(&VQ.J(#LJX83?[OZ63(JfMED]0a
36e-e;V,dE]XFF7#dUE8Z.@2Uead&FW6g)2FcfY8f@4J&3MU@#Mbc<F(14FgCVc=
/K2#.EY3K:34K:H.&HKTT=@CaDF+]@8WOYFAFRaQ5G3_^OX^O2LF>O4-HG;Z@LaH
@W,92#=D-b=5Qf(AVD6.A02<X)XV2aO0\HXgFB/.6Z0[AGg4W5FY3#;[8+?fcX&b
1V^U3EWVXD?,/W@\cH?DcO#7.QW(G#\d7@XNccJ6F=??(Sd1#aAI#,G[AFZU+UV:
=NKZD-I7A&/.JAV09/J+;XgAF(e7TU(JZ(^f.FABZX1g_.)T-#OQOS^K?c5Z<8[+
bZ@-O5eEYI2MD@aSJ)[/@?GE?E=FN[YbWG\&HUK#+?c-&<d;ON;0].f#85;c7Tc4
G(aB(25]7dEVc8U=LdMe?@O\.N;f7fK4;bS-,NAdT54J7HeZ27MeU6fN99XU[:e#
(U#+Yc(33N=E+)G/A=Waa7K8+5HD+N-KE-8U=1?JO00,NTG)T>TFSa[&e+_]-U;R
P5PV@#(;03W0GEV>B/Q@1\&[)BG^R/NO]#AF,G=8GP#(XN<H\9N4W5N@^Df[,6EY
>D6XgV/YSQZ@fU#GK^Uf.a8gNR092/+OKEAcO23_OR2&Jf9]A#YXW.9K)PLcXE8X
^K;3M(7F5YM#_BDfc.>P(,OF\M.0@RHcQ3H9TVa-OV<.2L<f]-]\B]3E)XRWYfV,
88Q)^J/\eF8:CJXQD>Fb_cTEGcCHMI=6X6F&)DRORM6<]O?#WWaA/0914Pc^AWVe
P3BegXYc/E;TP+?UAU><7,GI^@@gYE?4&[QDe;:7>-M\HE6V<[I+e@FDDb4=.S3e
YSMXJ=U]^)N6f#CH7[7U)YPg/5<S7ZAGbHW(N1^+2-bgYW<MZWG=O:93:-De),=_
(.3[&]=\.D+W7fF1[DBM@2U_g\f;,SZQBdBP(<f0Fa@;RY1M\JV<[QX);4U]&W98
EKS&d[]42PA>BQ_&2;AeLIBNVNA@?;VB#5&_W<-?Y[)._6)^eA9NcJY05<fRbQXB
I8cXf1)\ZB\A448>/Vg:SLU=GI5,CH_<I^2.e#c+D&[^S&/3?WBcJQD)OY.=@5(6
)<7a&:#F;79^GUge:Q<g@.^9R#C[+[5,=Y3O)><,QeJDQZ7E&_&NR,UdQW,C_MVN
NXK7X-K,RD6GFVP_ZbgXM&-):g[+Wa;/G#O9?I+RPbZWA=SbJ7Uf-1/a[eDJ6\>_
6F@J2MS/PMSf&6.\Y6IT-)Kd[U@I,b)WWgAQH#c</JeGeV:.aZWbcc(<6[:+2EH-
UXbES,DYB-/P9e><XX33=1.b^32=Ve^(/#,[L?8_Oe[UQ=B=[S=6I#GfNE0J39,0
[,BBYZBMTNDS8>PgHI<P)RbAQJWCR,H6WEH9&;(@1@aIANF82XTR\95b36Z<+W(]
6cYM;bC]<3+>c-?/K.KD4PR5:&3X5-8V5Zd@>cg&>P0YS6L44Y=[>U6POgNb/e++
93(LR,S11K=FAD+YT\1=NN\EDO?YW;&)(UN,E8TL?,B5EN45g(>df<eOc_:J863d
93A.X_]^=[X,S(_K&\-RRF;D+RK#PP2V7&]<bNPE0=P?Q)VdQa6-8BUQ#D95^=7C
53XZc<,@Hd;7UfFS(1--WFH&?3=eRV<C:596F1YYQN+a7N_F93cXCEbV/?_YB(4B
aXMN9O1B&\?-L2@c0UYgFZUYBZ^S0@&MCa@@)0AeKg=+J=ZS?[XNbP05Y:D=CVa:
:gNf0_9#Cb@_eKP8UbE,ZaO:I,WBX+Sb.?U=&@1g?FH2FJ7([J/\2ILK4+Q=2QEF
.QKF5UZf/:XF]6Z3M.]a6&5PQW.c.K@&8B^YJS<_7/ge1_=B(dfQ35d+M^6a:2IH
V3HT@JeN7#-Xea5>e7[(RX:3DNKScRSO,5S0^8I5#Af1fU-f>I2&+a-6=Q(5#B>?
/YA1LS\1.I.T,ODEL[X96ZA_H=Ag>,?0a7fA;>>NCFHMQLH[8-<4aKU2#5/+CJ#3
8fVaY))DdN1<XQ/d#N_-FV-1>_bce9_)KZ@29]PSHIW..>gZS9RcS,6:2a\eEBXP
OZU4d)V^aK&&H3>26D_0Zg4&M-(;=6;5J^I:5NT.OZIFf9K+V0]<.J5]6_N-,-/J
ERR7\^GZ#9E440;ZK)+YX(]YB_#<[g1dQ_ZP+7>;^\O])dINR;@82f?:#&+:96F?
CDRX#JXGI7bKARVI.1b5.K[&aF^IPEJQ7;,)/LeQaf8LQ)U-@Aa_V4ATKW^DYf>0
-P05+e3\ND1bgH_J0Z^P2F@)MSHSX)+fE6J+/:gXPGTKU6<3#:cb@MXRU63a>+>/
?GG[faB568H\eO@@^ETQcd)@g1gX\\MF;9.M(:839#L:98E8GBZdVKM4RA3;)1R.
b3g]9[&_5.@U,V+FXKAOa-G;DJG\1aZIBZC@Pa-BZ:O1DXCFP&dAO2BRZPTgR/QQ
]EfNT?Y]R>PccZYe.+,2MM#G##[#9S#[M#4:/,SA<gfA\79fE0R)JR0FLC3U&L.f
c<19F=Ad(+]QUc0_,#@S[DG]#5KG\&,]0@QF7bb3XOY0dT1T@R\#XL.[CZVd2S7B
1gGJD920HLT46\W;Kg@_791&UX>^c&L6342XJbH[)SY2D0Ud<R.;A_WN#fDTS)4;
^gWPJ99LKVH0B9KO5@NIT0/O>1D#?bP2SDRS.@?97IHDV9Z+QM;?A4[K<6:UPS;2
@db#<AUVE>17[3XdMKEIaf]MeQ35+Q@gR]RN&S/.\4];=D/Y=T/aB/Sfe(Y4ZRT\
WV5+1<ZSSeKNT)#QMR^MDI#fJK_,UU4]>C1&HI35SX8(YY0<CBMT<e7HQ67?2gd&
9N7D##S)MYV0E?O.D5DN8+H6H&H=/=edJCI#T+eS#_d05;FXQ<8X0gH&:&X^e)+.
BG.?b8be681^_#[4Z\f[<5b4K,1+9O8B9)<QPg9Y)+,T]c7A/AYKDXgc?ZRRd@^0
5=T]caWVU;J0d3GN)e&FM@149-WE.>>+^>V#5e[]G\;9(.=NQHUK^XBZVWKPU=:T
5,;R@I?7XKOGBUAd)R/-#ED<C5g<PeKXL:I&\Q]g>&;e41[G].^1K_,82/&We\[V
Af&RPINTUC/6:H:>FWAW<;W#fFa^SU2YO;ANR1RBe15RUaGA8]]F-6P\Ka?e=/Y=
0C5)>-Ub/d^UedgWR05\,Z/J0JG0:&42a3IA_V^B\M=C@M&3F8G&3JPG4TE[_W65
@dQc83cGBaBWeEP_EL@BJ3Y];?)/+61W>E,,<dL^Q1g5K[^g\C<S)eX[OefdC=3e
)7CPcUTH,5I8C,\=H2XB1\>Te00bU-@8Oe,29?GZ):MJYJ\5YP8(aRdWF,&/gbH@
(7OF#gQ)cPT?fb(cg,3E-(8_g_eAC#6HHgIVP2;]IU#=[6/6JI=\()E-?KW\6_g/
\98H.aMf8X7+;O_-8-V9bC-^&S@=L8.:O@[#&Q3WO/f9^AQ/&c)=#YLY<Z(?1b2;
7AEBRD3=,0A&8(:,YXBC8B9_MGP>;=6VS#H5(7HM)Bf\SV<@E;CbC?]D;WIIUH+b
:A9,/aD3W7F,1]>T@(LJGb].d>+#UFLf83J-&(<<0@^Ab5Z\2E/2&(ZM?<W;2DB?
aVf>P0/2^F1GCQ8)g;.;OZ1<TW/_)b5:_=g4,OcD@:]&)3YXHL=UUV8@5:cgQC53
-SN1G2]DJM^fP>1X[XR6g:IQS2GOEfAD0#e1V[HY8=ObPYC1,9XbWO;d7=(J]7SP
^8UX[B.Z_C,M8YX(dSeV>BLaD<?R<L]KQ@RH[+IIBbZCJ^+EBf/,).(QSFQgeTbE
^+WgXL<[.TUa8R@3_)3&6S4a=DJ\O;dYe-#-fS?c[0-_-IE:<_L,HY5_-+4/O^=G
Qd(,>LRg_E#;;d7H+_50+.AY#UNPaab_([c\].8^;W9aN4a#WHJP==BO.+2dR8UX
L-gGJcE,7:F/Db[+A^)<L@+@8T6HL0#1A_FKTEH0+M;NQ4Q76F(-/Yg8#L<ePW7d
;LgadHG?T8_?dDJ]7V=eY&cHX>[6c[\2Gf]LMYD?D?FFcgM[@b?48OTO\_;dKL>X
.X7L8XO8a/;Q/?+D9OC2C<P()W-\SI81+9g1DK0+H@&C/_0TSE<X]IS-7=_ZS+1#
OY=dE+,IKUCb^8([RWObF5NUc0eaef@#U9?a77W32HORg]=;a9D>Qg2QZ?<@#JSE
\a:.-Ze,;f29#VA+LBCG7[5IN:>gf66-A?UU7DILG0>:,=TM@#U\5TUAA:FfYN2&
.DY^NR]6K+)<H(gK(05HePMI\?^0b,JPZ@2S@c+.I2^@9&Z/IY\TQ]SN5d\:P<ZW
=.AX1&gGd#7PdHNS7R@D4ZeB25TT-+MSWK(@Bac1;6fI9&:X1MG2L9DE5EV+A/O5
ZdO,]\E>PgM(7TcCGb]b.)U.@##Q+aNXZ0@B^aZgS2cO)GH?#_LU;AE1YY</gBW_
>T\XRGJGb69[=QXNA-2-a2AGNGV0,^FffCZ8g<HU7fc?1P(4eHH6/VCf/[HF)@0W
AB;),?f(DC0,AD35;)>0I.+P9.d#Y824[LgH.)-c?E?M4I0e=#74HTXJ^]19M,Gf
7ABXR9OS.Y\TO+G4NPB<dTI9;BG#f6Cb=aSECa<X]S)5YRZ7OE#IL?4b\-Kb\=02
SS2YCbc8=6>_2W,#J\]/IK4(M9#?<<d^5@,=7QX^IF/5E]+_5=#VZA:=[[=<GW;e
1#IQG^N+UR)Z,;/W6#T>O)K^2EZ6TCOF3f[a<]:#14cLNC/Q3+b])&:;XZUM\I6U
?#22Qdg+S8WCgBJceVX@W/5J/:&Xb[S]),)]4C(HLXR[SI7\RWU]0E5H:f5VL\J)
0:bF1QGG(;dfL:_I6DFA\_T^_@)8X[.5^cYYgDbIVK_&2<+XT2,JD8Y)@3+(60d5
/@?U.XRS80)KWgLYDe<BeNIC@6,7J_G)e<HFaWTgd<@U1dKPTG[&2J(=WA75/3H[
+e18fSEJ(D=eAMBRSR8Mb[4\2I<<#RQH[9Q[Q.9?P/(?+TSX<>P@P2IJcJO]U8CI
Ub[BO^f[Q6QQ[AS&=H,5b+TX=e6I2GO9]OYDB^b9_/U(#.Ta;6Eb-g0RGP24>L#f
-1]TSDe=BUg8XDS+Ggg9Jb;HKe(BeU.-3)AF9R9gDPQC3XVGeVK63QJ;U@6_Ka,K
HBXW\Z_I9,]0KP_NW:12WC9G^<YQ>Z@H,^<d&,LCaMW67-\PgY4:AVZ)E=A^3VX[
XecL-5YLKa-^g-5a=,IZ^DcA^7Bb8cHUUg.XAO_?KH0-<_+Z4N3bAK&@?K(>a?E5
R-0?TH9V=XTD3S4(aTX?LF^9\^Zf30/6Pc04e7IANPN;\R1Gd_Ld&YIC5-EMMFc7
C<PUMeLbN)0eN.d]dbT,B(bVda(BSM^Ab?Ua5>,F=68gc?1N72MT]d-Z)_#a:X&=
W@Yf\E+8/.\QdEH.&2_cU266?B7dMR#Q#&S:,=1D1<Z?f;Wa@S+^5>/YP;=D(9YE
+_A#@3^9^?5P7M3QQ<Q9<=9d=?)(aNcQ?Of)3\If<[<<I(PbF<B7.&+g+8ed&B]a
Tf2-Q.3]_6;.[-4Z,M2\ZTO\D,4?WV0fY<EUQT-::caD6SgHfS0+JX//P>SAV\&G
RDLaONO8-Dd=R<=Dg3VbGI_Rc4>4MRdVbU5B^?@PWgJW?9aR4T@./^/ABH[\Rg?B
cUa/3AY04cAZ;YD:1C\Rb8#X>HA2)Q5HCXL(.DBdbcD2P:8<R2_2.+6c>D-5?\##
(DO?e<KcfFQfX+MRYc+&DU^Z89gB9/S/BZG&TMF4f9gYgR37UO6&PR1H1SC)7O_X
J;F>>6c12/0[3ZWZPPV/[R8_^c[^:0T.[@WPY[HSE.)8OQY&;V)X26EJRZ#>@#.Q
b/O@POWC.&+a./PMgaO22L9:8b&W1]Z;OH:DA0>cOTA[J&1^HJG@F0/I^-dXJ@(V
aPT)gCde>XNMXZL0AgfJ1N6[4ZgBY2;##_TGZDg&_F@^:.:209g:G&3BYMA4Z1Tc
J&=3[,T?:.c(I\-S).E[JK#[3Y4MLCA^2e.,TIf\cG4:KJg06@,7L[dL5K#J.7-#
E2LM01Z0EC;W-0K1S<4@V;LCHPN6f[P_IHQ9ecSE1>W^a,_;#a3=LAb::XP0)S;S
H0>c?B@TBK[_C^_ZY0N;I4OJ&6M?Wb;5>H,IGRORbc]637b-;N=F]\NRYYPWe3^:
>G]1R4:4S]VSeK:1:c;SB&d&>@?M(^4KS[^,7<JD2OEHP#aF8ZdN21<D-7^U4]:U
KgeSX.P:4[BQ+Zd--3OZ&\W)#QOW5UTA^3LEM5FL,#++J6HKA<6:9?=I<\5=60D-
e,_>F@/+5R,F;;/EI?CTHb\K#e50GRBA9E()5Gf(7KGVE2\E7/)[J?>(SZ3^U@7P
5@2+?YY:[f3R:gV6S>DZR)0QW:\>Pa2gJcGaPGEVJ@5ccP=0UD?\;OSbfC--;P+?
1Q_,EF(N5PE;G)9+)T-R@@GJO>.:,#.g]3Y2Jg<AAe.G8^<JLOK35gN^Ke8g&YK[
&X\8J.ae<VWJ)S>0^B;RWb;_J4M&Y]/QcRC6IOA5J-VMd[20R.9@__gD=X:X?QLG
-O3<1I+5@e2W2Y2DB/]G-;J?H9+f1K_ZD#Q>,>)#\EHJ4B40&]J1<\54\VaLMX7b
Ke?(c5SNgZ#NJ#200VIf=,HK(;+\&IeGQ,b^9MIaDV)c;)&06?49BDN8K<+-N8M3
8>ba(_2:Z)^]<6bHK9:>d)4K^F?)2Gg;DF594H7UTS]6:VY6LV(TKRLb07HVJL\=
cG#Q>.U&/O1N#GG33;#CcKd?8?H:<3Z##eRP,Sb/^1+QXYZJ)SN^GI.Hg=.#H4O(
-U.OH?[#\7OcR0-^09S<<T;K3Oa3QD6\0EJ3a-K9#:H(8<R[^1F7A7;aaM:S@B.d
a0_g8#(;807H(X<gXW:EGJUXdA,?aSC&Z-L+AV>&?G.8A65+_#K]\g@f7)BN,NO7
eSgf.F9]eL+OaA?P#;Cb5#?_3;f)beD^M,?@(Y7bK,RdQ:A;aeV_(a(PaOK;ZM)(
SfZEcPbHa6AP)Y5@.VeP>R04?T[>bH-XCYZ^WC49R>^DaJ[\]9_MaX#YWHSB[SY(
K06GdLEQa2-AaF[G:dH(d@HLUH67Y.M=cRI_#(gLU:,#<Q7_bX&N)=T2Q.RR/T]:
B^FZ86D:@]=EcK)#CDOLX<ZeT@RFb?SA:]U44;NCSJEO(FML=V=;H#?B,Db/<bEB
^G:X.NSG8B->c:[&DNaU<+S<Vd_^HfPcGb.&6D8Cf&abQ>PD7f/aQDS8baL0=.If
:7(QdXP@+9.@]B?38Q.PPX>a8RFFf&^4ecFD^B2E0EeE3P=;J.^K#VIH:6<2L5>J
MG3:Xg]#^0;RL[TSEg:g\ZM=>U0_SIF>H:]=4g;0.+@-#5Vg-;JDD8dZ)gef66c7
S?]OH+\);HY=6;F/P?(WeU9&8N-I_d=(7)a/>=PXT:T<-8O#XRV5OZ5#>-A<H<(2
I.4C0K,(e@/fb/B>_B+J8T8,2aG/VJZTF;^&-EBQ>QPW9T6Ef(fK1g/6G80d/R=2
=P@1(.72TLd2L:SH&@:>TD.-6EHXK6RMfbV=[G^^_QNS4+RaRPg^&;4QOaT+Q=U9
RZ64C8WF6B?TE\;60DDW-2DQVd\GaFZ<Vd]aM_f#P]d)dIK@BMC?CUcHT44\(3Db
c074WCWP-[22CQ2DWe+d/#\?Rb=dFR(Y90(#4.g[A.H6/P/a?c;?-Y<-/<(]&V3I
XZH@.+(7YdNOGK#TQZT>&;]a<4ec0Pf&#c.(J32=[TVA2?C7BQ,])9ZbO4<.AH(8
=J5C8PX1X)e+,1TY\N#,_)1bHEb(R,]D,Y^Q:09OORX3d>O:-I.M63>O[QefNCYg
fE&#B1MMZO4><_DP&IRDK-K&cU]\:P#PT:?Qg[fSY(FVE2?@Ecg[UHD\QCLeNd?D
_(?PCb?]2KS/8]MZW#Ig@\4K2-VfEZ#Ia]G;a5/)9ABX7&W]O(Y]=0^CZ<X49]25
fJgd+FN]6L\^d7SKA6QX7bE)0g5Kd?V4B:?.\89_NES=/B<_Y/T99-8C(\b>?&V5
]1I8PVG-&3;(^<R8N?7MBA0\7f?UO^)6R/4\<((PdKBS]Z?B16EBgCW@feLOF/>[
]T?GI^#V8[?]4,1=>TRI3a6=[SS5Eb@g\7]bROcYd.6DW9TWfa;)W3>9Y>#PBU^c
=9O85@B+>/ea-;Y=2,dAf)UNDIV(,f1&NF_L.CcP0?-Xc2QBY3Q\e/WN10eOCIbJ
&G:,H>Zb.M/S93K&d3Gb@?8b;=7+/BC2=[2AWJMbJ]->^_^\,MLe\I6#I2<cg[41
\5,07&G]R)AVTJfC(_P1?Xd1FYVCb;UOQI+DCeE0>N<Ned&G^F9NW:PV+\Ag9NfV
1eKgP@[[:CHV#V84VHF,Z/2N16XN55HS0J)(aC#&<Z6=T>5+])QXL3SI#A)IW_W>
5fSCE;K8aO1=TGCA+WXL@WQbbgNEE<&1:gcS=f6RT&:Z;GMa&Z2H+UGKVM.1<Kd;
a<:KTb?D?9E+576;H-=NT>#e7(ZXX6YS9g2(V[)8e6)D@QY)>_U;M3U;BF;+H-.\
0TQ>GN7&caa8RY0bY.Oa37b@Xb:bAWJXOD@23^aFP]0=6FNJcXIQ^ZOGCPK&2-C1
K[4&S^7^&9O6:1_R@CAK.FfM:^<5\MY5ONM@D-P.J]UGV+Y(^]Y0/F<4H-W.L<:c
AcTFYD2?Je)1N)D:>E)6@P3GK7_8V^U5bCJIF5B<K0>1#;\d:]f<Q0bHT#4]T=6R
N83bF4H##&M&FgG2DEJD99Z]Yc+;Y2Q<cJV-:.))#IK>B_PGNQ.B^KH\V?Ra..R>
@ZV?eI7d5=P:OMW7+.U=:RV>(G,_<O13SRW]f:dCI@B7Bb+;C+5aBN=O#,PQO[A[
:b.P;6ce\\c_2dQ(3DT3-WVfN9/4K<@=g;W:ZZDW,0(139@e/23JCKVH9/LE;(O(
JcI]3&bf&V?g0fV>UbAH5+S+WW@A)ZA+HVOO24WHcK17a?dHc[c,A_:GJSMO4.g/
PNXO^+_^RS?;Pb6GJ?M:5NPb7.RR>Z/@.B:c9SX4?0f\7N^]eRg4B&2DDTbBg-U[
7U\9d#7)HM4?cJa?5Z((fQaKVg)C2)1Ee11\6gP8@bT?(#O/H<O1?D)#KH.3VOYP
OL^bA(19R/Tf?PebV76<48K+/_^dbbP\27NV>FC#4(@?cRRDg\U&S65)[0G:UR9Q
1PV(eO&7@=1Q?V6DF\=V5)O&LC91#2_aM0PV&00BDf>-[@eA^1a=YWONW#=NX[&c
g:3C56SbfNN,&AB/0#]\gE-II8CaT+PLO_6OSWe<gc<c_+YE,,,.b9=F#[3OZTI2
GZQ4@(f2:D>\))bcbKCKU^?VFX^)^W0:dfeaZKT]H\gd/4b5;,>G]CRN=0RF+6Jc
F@2]E]XVO)6#8FM4T-(JZ^F:QB_P]&;<bY-LJ.8Y/[)4Q[D\3--3LWOU+]#&TT\_
7?::?IU\ZA.H2Pfd:D1:KM/3\WIKGfB@Pg_c\KS2_Qe[eRbB)R@::KTIVS)#ae?\
1M_W[B]N2\@;.V.PM7f1TY7-A,0(0[_VIXOUJ4e7Yc)_M7WY^gNZ]S)6H)ZL-ga)
Kg^ZYL7D#CNZ8ceLCfAYH5>ZbSSS9-1V&L(]PA2&N]W7]V4/M;P=:S_(+1.C3RN_
EJUMg>WR\PU[WA<PN?;c(fgdS4LU/D?@3^f4NQ_dBHc8</]77X9Oe6SY2U;E./&Y
9QgfGI(YP+&<07425cJUeBRM,YYMUF&dT2Q31ef]G]fP>2^D3b&>S62bc=&:\?K^
9G7\0d+_M)@><_O=1/1C8>U-5P>UN:^+1MM\&(IUS20LHW(3K.-G8DDS#C@@C6YG
bFe?&]@0@-IgG86X/#6@-GI;(GTfd<<=@UGOeHF[.Rc1,A40_8bZfUNEOK3KV@@3
EC,B<PCeSZODK,6H\7-1T)900PSLL\>]0#)B.6f;UIQT]DSOP^bD?))Qf3=_1.?V
&KEf4>_,WR6-gSDK0Vce7d4#/\ZXdDC05S-JaKeIW))Z1LK:f0E&5KF1\YSKR/1=
:ETd:UCII0MgD.6+KZ<?G/6LI,,XP)SWacMSfIFY0Xd8ODe5g/VXPR^bE>S)ZZ#:
=,HS>O1-67YGHJd_RHAP[=C,,Q7H:O>CA4DbL>1J<-VI:2S6L#gCT@HN=[c1L.?S
+3Bf=^S\E(V>-L;/5;?1C(PbU2]1QTGP-dKP?U)cc<XZ^d84(:=S;P2TC;F4g/C4
g0R6F>^P@G=J=C-E:\\FG>UL@7;C.7Ae)L7.5:/@NPV9_.dVV3geTO)?PJ91YUZ.
B)RBS5@M-aLH&4U^&fG4#UK&MV^Z>UR:U<ZF8fOdA3=RHX^_&XVWTU0Zf,A,COO0
W3YV>K^ON/JJTK.X[8U+PeQXFO,>RZ5(fF//?@VIK4@Sg.7T5(MMCQTfFB2H2gC&
Ng;\.d?Dc^cDQRffA?Wa_\ScV>5LOa@7fF+A:Z:bbVY7X1#LcID^_Q-/gZ0H+]Q6
XN6OY]RZY+N4LcC:IMEAZ]X96<QQQ4KC@X,4@3=2P.06cd]EU>.[TEfUN2ceAO>Z
gI.#aK7<5.06=)FX9,)>AI:/Q:OI@f4U<GADLZ-]@BdC#df<c(L,:4C:Gd&Pe4=0
Gc[^eKMe<-=<;&=)7IZC1#,=2b[ETD]IW8I\H&dG[U\HP_98T7K;ac9QL\d7bL8J
>9cC>\=\;f7bOV[[AAL0:9b^/>/^@g-T#?_;9g^=PYU06(J83>U68H;7.D]/1Fg3
1NL)JUAGaYXDQ#;==.BIcLc;/J/Jed=N<FJ_:W<c-eGg\5RWaT\RVN3^d@>KZb-.
:GX^7+?YU^a8\8AdOP4)LdON0AZKQV(M2LeJH<RF9OD&JCE:47MYWfaX1>STKTJ]
P8\>YK3KZN5V+WB,819JTW^LS=9L_b-O8GCc4D?U^-B+:7O^LUTWP8+50+9FcNKI
:X;NNXN40XA6c;+)]:#;#RYC=CN;1IB_9MI6R]NFR28@dN[RKL(FC5^e4F[YC?71
ARR1D<a289f;TS82[<]AbAK)G7U;_gA)/_[NZRVEP<?2BH#:ScT#9Rf?\<9XbUNS
0R;+C=H=6bT8))0=P.C+HFg5^MTYT]AJG\DTL&RDMa(A2e\SaWM16/=V[g-[[PbW
U^CSVNcG)B9()^4=8U:S(_T-J@V(TC26Vf-RbVU?V_c7Ac8F^-ZEQ2Lb8E]&,)TY
&OcVB)X7;#gWRMGZEaSO48;=DV+C5,JP@)c/^0++J/U#g7\Cb=A,N;V<PMEQ2d2<
Q0A\6V/+NfW;8_,?.YJ+cP(<3<N[U(\Tg4V0?6GbMMT8.QA/\CP?LO9FWO39<Je;
N53LETeBXUIa0HXRf,AKXfc=g;5<H\[J26Y&ZW1R(B8IX7fEg&aL2fK[cb@a7^@2
gNYRMGf12/H1b]8/K^S/WbP,L:f&Pa8VU#J/Y#GbAdT)g#NX?,8g;N.[_33Y3,?+
eZ>;G<JHg^=GA]+_/)&.PEF5@a;:L2&fC>P97C[_RZgAWTC@\//[L3ZNSP2_8ERM
JTU^6:U_aPC=#KFZ]TKfMR(K6\S56[^eQV67<EG-a12K::?f2eUI18Id\JNb^ELg
3&T+R6OQCPS(U+YAYe,91V>WYXdDd1W59g7O5OLH_EZ(/bg#8@@gBZ6@Eb3N30;1
J)F@&&b/,&/EI=Y@5;XL,482d?+2gUgZ:5NFSX@/.\6b9P05Je=gL3@,Q,3-D=_M
ZC@ON4C,<3+O[MQ.3(]6G^F98K/2GZST2U=YJA4Y@>fAO>,)_G^,SL@8Q/8/2T7#
8Jg+c2+R-1YVGPXP:W_C08EgA29GV]IbfFFM0BI\(@6-8D2.6)R64&-gOcUS>9VU
,#BfEe2_>058NKd9VNA30(B;3cZ1V,2OgA_8\a@3&A3^#.\-If&(3?:#EWLT5L+U
6SU,GQ9]_6[CS[K#[cTPOgQ^NMdY3N[.W082Z:V/UUP\)c\4(^P_8SBf<R9B1WdV
;_FPFQ/M.7BCKS+J<>Z)FA5Ad3&?2R5>ISM#U/:DB[W4?@2-_/8<U_O>UU1V1e\Q
MDZ97.Y>Yc53&\EWGKSAL5ODIgRM;?2a&@f4P3ALbT2]5F-J=C-:[Zd^SPV.XUb2
]FT(M\?ZA,?Nd2-AB+O4927FVYQ1-1/]g@C8649AY75gKEg71\cda)97e,HROPUG
Lc@WNb.<\2T#bbX/OOC.#]-dff6];3a22LgQ+Fa[[JBK_2ITRA+TQJFJEQ/=R:=&
_X25QFHDVPg?U[C&T/5F1GSZ9eW@APSPB6L<AG=DZ:F6d-DcVH2AYOR=EN?P505B
A0]fZQW#CTFVc0AX+[,2f&#]R0CfZ526^O(ff/VGK/98P1.RT8Oe9e7O5)?KG\6T
cR4K,W,+P:8TJe,>J56_]2.AXgY;V+G#b_/d:J87cGbPXXX@_aU57a^P[QOCIAS1
W0C^&+9]GU=ABW;(UN@c)O=B/ZAe82Ub2HO;7SUZDT->(.Z;C4TX/b:JR.=XS/.\
6,c(.<ccI;QOCYAbaU435Bc:UV^,H3L<-MS\cb(aUb1NO9W?Y0-I2a?>,Eb8>YAX
JN2_[2B>dWYeP7;64UFbU8\bdfG&-]eFNZE7bZERXgATY8Y[6JISK&F9HGR>TC<_
U6<U3ag0_F;_2SILDVHI-8:^Ua,2#9ITSU2cfUJ=@69<H(MecJ@<24=<Ra@-51:D
.S;b(M0fT&Qg,eX9Q9O5YD[8fYM=?W^NISRbF=+:05,2GKVB2:<28DCVQ(Z/a\[_
>9O7&ZZgE<:<1?+PgKBL58N]<W](2\(3UgcM9]-#I]_#60BbV]SR2LZ+Oc6,]PFF
]F;M+JZ[.aL03gMKO]=E&?RQK42#HAKR[MF/MKMKVTG\dc(=\9#cC0118G=@BV)6
0[Sg.]Q>F6Yb5NGQY8H55J:QVbYbe>+CC:IAb5O]DV3]5T<?:g7bS1f@Z75T-.@=
B@60>cT-+:OR0@::E&O^.,9>:=HD58b68_(>^U?]@#5&9=0)(5HH#/NM[>\Q6UKR
/:/Of1TE+?,I(McIBLaN8?97aC+Ad^b/W6_N#L64#G/N966LBfH(-&<6Y=+K(Ifb
BFF_8D#11/DG?bOW58Y+XW^G?LfJJ,[O;GFYCg:BP7^0/G[0AfQ:33G\TT=]V@]a
06UaT)DY]U)5:.6eZ7<G^7Z+\<,D>F9C@&_Y-fT2X]:_-gOZEL\#>c;_#7fT7.<X
&=C1G4/OXE3a8W;e<H-F.EJbXVMJ2cSDTROEGgJF[5/J&1B(NA3O+,bVf&N:[)=B
,,a.36Pa=d@,FVWe?0,P^/9F2[=SJ;G5b\-+NA;TeC64V[65KM8)2#JE,V#76]&N
@822-UW9[-^:?SK63B[DUZS>^ANU_0AQ@RJ3Z8DG7#@Jc)e2B]c#;6^J[V1>8J5c
G/^e<dgW24\ePg:I+^45O(L3D#bWORSde8A(0(,DEfE0Cd#ZH=7,XG=/CKZV>gG6
55fLbBH^9W86+46DXK0b8ZJ[B#(S=BadSYZ,H#@/O]XK<P^VE/Tf\HE6CdE8-?#M
1MIZ)<-cXLJO/\2F.HDN-M)X@fHWH-H7/:0@<UG(12C)HQfGN5[P[TeHG<EUF,(F
VPBK>-\GVDHF,OW>>g?@8_8YX>543-9bXVYIRYFNT]4]CTL]O45Q:OOI,=A4D-gb
/agEI<2HH:A(#LMACa@;[gggUgN1_(_+,]&,8S9KAUBT\N:DPR+Ab7M)K(]V.=-8
K+[W_Pdgf=-5DPPAM>7OEJJ0FJ_(K5RK>,HR;JB,5?RBK.J5JaaN^:XRUTXdE_PP
4FAccePX)@\]BOLg2QT&9:K>04SW14E3P=X/9OKI&_(@8He/?(0\Z>ZSGeY(FfUE
cDLJaZVcSTM\7.J[a@Z,<B40@PEUTS.-TQa4(=0bJ_X+3[M4L8@4;6F0[3U-HZ?/
D=@5bbQ#ZT[KVF]?O0P/F>,bCFb<=;9[<2Lc\/PHJ1E2CVT8b7<b<_K;^74CUaX(
:@J/,]8DC<edgf,DPY-Ma18ab<@]5XZ487C)3B#9KUbaJb8INLYYZ^XPRK>X2C_;
WIfWRQ1&KSDObIO&^?8UDH,(d+68J[7HDX=2@KG_ZN&<JLUE#0PGQG;CIe-S-.?(
NK_:U/4;1G0GN]db(T;38BIbGUZ<La;)=/T)&L62918:]H(cMZ#KaXb,D=@C#9?M
I),&cLSXL7]OeF_.fcc+/YDJS9)Mb]YH?(@CX,Y<W357\3H>A7C<,I1K>=V]gA>5
_6H?/1Abe(QHC13.G3HXG\;eU/B96/?UQYK)C]XM,5IDCVWHWP\L<,bd=..[DW=^
KL#(^fBE?V3V,[M65ZB4f.PD0M./3KJbU;H+b3I)6d:KEAVO>>.51W(2.J--MW39
9.OM9[=H1YOg36O)02-,<g^<;9@-4<Mc@Y?-S]V,V03b[C]<;cPED@FK&]?7))=9
N,b6;U7^?G7:.YT&=41#5LL2/DK9:F4A0,IP)).7#+3@dJGBT3^]9+06F9Zdea6.
73_NN<d<--QYg.2cePf?PQZLAX7aS+94NHWGfX9<D^QEQ[)A5:]_DcD.Y7ddb]SP
QT+YVXE[&Za1.abAXL0Mg4P++1MX=<C.N?gXaR3d-SL@IbTQOFeD-_#eE,4U&YD=
UE_IcDMKL;8N>,26R]#7),a&.c.(EZXN1QF[bML(Z7F4)6)G+(f:ODdfA)5#J4DN
7B,)^C_<(FIC&AWd>=;S^=J;KBN75GC#@1.0fV)C.^54H^F3(S(P&(VGT.ABMBbA
>>IN8Q>IQg@&K+3?1GGP@74^FCOLKDS]d=;?fe?FMH<G]aC97EJ7B<_]J]OSEd(@
FR[Cb6?N-U-9#R(/3c<E-d3e0A3(?#,<S7PB\fC/D@.ESa>IM]5\Rgb;V:W&XBIN
>]&[CO86g+KHH1RVQJK\DgO+&dWQQEa6QL054/gaJ?C=@_)5@@+Zf;4d[a(VF)J.
dK^PW/IH5.HWHKeH9]ADUaDG#4?Z_KKO1#8,=8L&TaW+7B.Ka0E3N\PV:OS,\(NP
\0eH&f99BecN&POEXL59:0P,29/cB>Bg/HaJ-)_[42FWR#&AbJVM5[LRG6LZ>6/?
R4YK7(9@V_#RDZ)e;<+^.?YB3CY\58YcJ.<.be:FDP:,PY29UCG4E6JZa4ZFaU<C
M+\d_#Qa9QPL5IU9?W?36+-<??TT^M:7D+aTU.7E)Tc#Qc_@#f\\3f-4J\@2YI&M
NP3.c.0VgYVBYF.T_A6Yc&IK[)U52.KD<&g<I^@R(@1Y#:N6OS641#<H9gXX_fZ2
77Y/0XW^N^Eg=<C#(];-PW:,G/GA(A[cS71FN..K&I(,&9L@0(K-]f@b1308b<[c
])8T-#]b@ASYC0,.g&3.NF;JM)V?\ITZFY\Z/<<VY[#J5DAHK7_:GAbLFYX8#IOZ
.>N6MKHINN5-#V@=]W[3eOQg^?H)^LP2Sc8_QY7Jd^<g8(=;d.UgOV.RJe6^4@1Z
I-0/S<SXc.YEdL;N&0XX-Z8T@eBAX_Q&2?3#IWe\\_@F/-:1PK59ca8_2JGW.V6_
0@DS+\gI46ge^<JTG[[LI^SeL:d33);UE=18L/;A5T)4Yc,.M5?R;DKF/@IN86=/
24T/C3;K:,H1<_+?R<\O>R+R@FKUI&XZNS,8_KOCc,/6HT4T?@RBXCKR5g7OKJCJ
8OA@8fS_/78VV.d#=g#CeIGN#QJ:,B->UN.AOXAUeO7dZD?Z<Y2APP3+7eJ36P9/
7>LZJ4V.^aY@La[7UJK4LVWZ;^\V9@CZ[?X@&R+,O3F&)WP&(V3MYV6W(OMHQQdK
d3&#5AQ]b9MN3&&H567[VdR1f=F2YO7/PRUfa:Q4P^eAU_fJ^A9(TbC[##eW8A^/
YJQbY&P4DEN/5edJWaRKA)E\Q9G)YFaYVH?@O5K^F+FWEZVf,9.-L=E[7f1H()7-
_2NfTEWJ@W@\(D2I4[+I+7g_<S32SS-O/I.-YI/fE=bRg-d\G4BB>82TR\2[BMEE
-GR(M0BK5fX_5&<@OVKF]L?1J88)fGYcV-9K4]REO)Gc)2[c8U7/,WN^\YY(IDQM
[=bY(<bE4./O2>E/RYTKN17g1D@9@.:7BGP#DR>eM(3#@1cQKdcL97->)IeHYaG1
6E6f:@]F;(40EN;)C1A8TG..#/@+(g6KV5=5g>P1EM:9b4?Ua,3:\.0/A9B6(Ndd
C#Vf6]+HR&W4[17Nd>U=9./eI,D07W,Ba\TSWWHPgRY8AaV0.#VI=_4=gCO.^ggJ
UfK,::Y_UefO<MBLY=@B4ROY(,X9:L\cO-]R_XZ:T7QL[VHM@PJY[5PNeWa34=eX
;be]@^6SKY9AL,&(]LLHH,MGKefI@8ZN26DL?H]OXXAR/BIG<[Cf1\(Z,N,-gc:S
TZf3LSE9PN,D\\T7I-\XZKS+6&QY/Sa#==]gOZ:1Z)SRU=0&I>DX3:KAQBfXf=T+
R>.GVcQR6/G\_]@\c\H6@.DLF3TLUc?Q=cR49G^:+4@3bAQWKBM+\<a=Ed-LNX@@
_,YaPAY)>E[CXgP&O9?66H]U;EM,/83deNW_We<9(HgFNc+f2.Ab>gYC@9C<Dba7
e-11V.1?e)ABb63JBOQTFWRU/_9B;f+_<YY<[b-M]WYQ4C[S)=35<KB@Z/L6;>a-
2^@cP]K@D;_WJDGPE;4Hb<5B:,+b,Dcg_-DR2Y-1(1/#EQJ4aad:B4f)0PWD?\.9
EI)#eb<U+G#3YNF-/LgI+dFd7-,KX]G3+M)TCd\_TUY6=N^TRY?c[B0,-82^N9ag
9K+<KfX2V+-b9EGLDX]ATCU\[W\O.0;O5M,.Z.KI5T]S#)CSLA7&,-PY89JK-c=^
#KfF.Jc?=[aC(L3a[FUHU.Q??H)^Qge3PO^AW>+T@7R[.?ObR=dHL)-dFcFF>X-d
0fL<?VDOY8&I>V.I7.8PbJ2EK5>S2Qf&2YPO.J;/[5JVE@FR=>-GBTK=+,MOg1JI
@]WQIDR3R)=aJC8@@3)^fRBg=-#W0c&6X(QV.aBW[7S<\Tg+;aNU.TWIP2.J2@N:
@S[J+K53)K38aU#O_E/I[L5#9A9[)2@_@?B,eT#W=.^2@f21+\;,N=\8)]?OQIU4
0dd^2N:I\8R/Aag]cGaQQ5VQWba.)C6?+)?<A^/&OK+(O2-c=b5\]8MJ^dZAT7CS
M5(VVBY6La#+f2aWBRXW?b9[YKROOG3GIPGY141=1@&CcAPN^a+)J1?J0EER(AJB
OBYc+IV_7R(1-E;RB3@KcC3:<0E\=DUT9g?C:K6S@,VPPAUKS:NUNWeZO3G9R<gW
($
`endprotected
endmodule



