../02_SYN/Netlist/AFS_Wrapper.sv