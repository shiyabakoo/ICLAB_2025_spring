`ifdef RTL
    `define CYCLE_TIME 20.0
`endif
`ifdef GATE
    `define CYCLE_TIME 17.5
`endif

module PATTERN(
    // Output signals
    clk,
	rst_n,
	in_valid,
    in_syndrome, 
    // Input signals
    out_valid, 
	out_location
);


`protected
eUDV18D/_J/QE,EVa7V:eE\9DP1T.)a@#bZd\:>S]AW0MbKQ9K;01)/D4H=3YY[f
3AfDT.7MfGTZ\(I4RMOU\fd,\e:)070eC1PL_(Gfg(R_N=&(eP_VVTYaGVS1JBU:
;eg=ATQ#>@51T?,Ne047AZWMdX9WBBa1(3;+?B]T90\R^MQ.0J<+gWHd@_Ibcf)6
^B.Yd)2d^-9QaIWWQ]R]A>WM5$
`endprotected
output reg clk, rst_n, in_valid;
output reg [3:0] in_syndrome;

input out_valid;
input [3:0] out_location;


`protected
4\J+SAR1+JVYg)O.GT(dGbH=PRPA,QBGU,a\V7ROR4NIOZ0/:O417)HA\34A_/.#
[83X_ZT@,(P]<EKSXUMTA)E&#UE#8VbdK5J80BPF_=>g>,#-#;][>M><FNA+MKD<
cOe<,1+a:AXL5efaF<?/\FY.e1Ed\K>b7?BHc/N_-I<&V?11)baZ4=,@ff46?^(:
@FBX0]4f)7L4??[8gga7[ZY@a#aMbWeHOEP3DUE\[R;XW,O,5R?Ve(bc0\0,+2E3
+@CPff=@aF_SKA[TYRNNG:JPaDJaB5C&4Ccd0&fge7+Q<VCJ+)LEJ^5-PB@OGCO)
G,/I/N(#+:a0I3>E^1=]P>_HF7>EJAffb_\cT87g>)^1WC;CD1/\I/;R2a0??7/C
4MZ==a=LXS#C>6<)&IC,BaBBU6C,@XI327PVT(T#Y2(CM^Rg>,M>I[OIdXbH^Q-e
TW\bY)7](>]RVTUf\V[c(245f(2T&O/YKLVb^ZdRFQ:a8@,2K&:55:3)bU?QIS@^
+>GOL-G801+feD)S-#[6Mf45b+dV:E5BBAf9]O-RIbVacE-<0LQ<cULTM/<PJfM6
2dW.XH6ZV0e(8#3X<7?Qb-b/42bFD./N(S(:]?\3-9VcWK(b[PDTN4=UT5HP^JBH
(:;CYLB2ePK](J51+10(W6YGA@S,W#-C,gPf\?FF[bTg/44ggGIDUc?G;8TLPabc
:fa+V,F&C6K)+bF(]_X[HLS7SYGZ)Y1VH#PGa.O#0TU&-Ed<cG)>-(UVHSKY^Z0(
P.@CK_S-#>19Xa]<.+,AW;NN@Sbb&MKR]0-6gdGEF+EFX^Nc5bB?+&V;>GLWAFfO
32P4I8=H)DXN_]<-_QeaYecG]N<+<f3WT^H_YB&C6K:?.ZDIIg_XA)\db(O:L6_3
Y_OUJK\b9)f&F0?LeU-c;<,b+JME=\[1OI>_]X41TP@L#]J-DM4Y@^KCGaY=9<e&
BVUN1&UC4OYD4eQTH>R#;dDP&F<L3M_JW8,M2^@4IT/(/8[-ME4T2^cPEK8M>704
@;_&O/;c4Z&B[4bH+5V@8LEY>K1H/,=@\Q#\(bY?e=Q:?BgO>(]QF\c8T>:/U/ce
OB#1Q7A\(VTg+#YbOFEHF7-J1O#FL@R3,\[/U=^&9FWR</6J7/4&HA]V0ZMR^F^I
1g0.<CAY8SG/5D:H^3]WLZ12CHWMbP24@VX9:SRN:XN4>CDCdf(L]13-P^,/;7:P
Z56#1\?LOZ\U,0Y?NbJWA>G@6>CTQ>:F,T00;>_;I[ge3McL7AIR0-SXZ8RfUD+C
gX3?10JZKEeF[UVI9.+_#N72#357E0T&.1CS]W5.#GP2-Q#FXY08_A..0/2M5_07
W8&IS-62D?c#QS)1/=cQ2Tcg72PH.,VHK3-V3B/(NWRYZQN02Nbc[ESfZO__P-=6
.0c,)[E74f;L8RBTW@FZ6LO?J,ZB8CFT1O&40gPcX[+XSgVZMUJ4D/g&_DM^]&<8
EO5R#aB(=cKR]6H3gG)9G3FDQUD)RE7G;VJ-B82\,,e[<))_N\1\&A.WB^Y.b@b)
We;GLRM(?O6J13EJ&Z0X[Ma>0T/BgQKF+4BCfbVcJe9YJ[#e@Xf;PAOb#+1eU6TF
SD#9S+XR64-&0A0LQ>XCGH-;OWbd=75^PZb[e5>WT,.)?D9T&ga11[31-10aG>Q2
P1<GaF+]4K;NXFSKK:2/UC4.W\eW.ga)Se2+2?K/RCA)L+e-7RJ0F>8.d(#_MBQW
:P\B.a@H/,>#K0^\/MVA0,V^K4:98TE5b@\4[SB[aE5&T#cXHEdZdM=VGM#7?<>U
4)EO;^MG4TW>?YA70#Te\WUegU_<[,&#1fFZ3Q(P<><YPQ<1B<,H43X-2P/dZ#)-
-RY(;2E3^.CSW&b/;\8cAc-IQTZN21(8#XIOT?EK.W\DP<\55HCfD7bZKAWTGXE(
f5cSF5LFOF;70eWX1W91[K_gZOcS<I.J_QFFVI?\c&H,Fb2a5T2aZY6;&\A2G5GI
K-7NZ/@IT5>\C]&[..:/7?7[,#N0BS:a466UK.G,C3R2bW&JMQgT^3K&#D]F=(:<
B_<MgI5<FB/dHY_OLX+eP4L6-O,?92N_-15b^I+a8-Qe=cE(C6:H7RH4AeeX<^/K
=Y5Q(,\KBGP:/[/3:4_4S6U[2CW/<Y@AadMBE#=g]Cd:,eQV<M_VKW3L8->Z7WG@
U#P0J5Tg&LWcVab&84&2(5^1=8ffFOGS^^M9DE.Y=E=;Wbd;=CJ8=[5aQbO?X^<e
b>\IO73W=Y:6.d^6<3(c.cAb>7M9C4Y^F(@B<UI0Q\UJR\8;a@:cC_Ve4N&d/(GI
4ISCfD=NM#>)7^?31g[(<VS[EH6?X)E_[_]X8HOV2>df]9Lg>c9IU-B=L>>J1A[S
Na6EJd6D,ZT9C.+MYeCZLOYXDA?R(/VN&L1VQXL+F\SHQ6b/EB6/0]3^0#5A@5PV
<DE4gV^F_JNJ[6)Kc<;(Pa\-Of#<MUdE@\5(CS@M_VS1&ZP#QAK-bWK-)KELT\g^
\/(VgQH-?fbPAY=+Kd3+B.?V=]/56,6MQS2#[DD^dX>T?0-<F3F1UcgSUXeR:)6b
c#>>[_RPU<B4C#.;50cVRU39,E[E??(/K1&eD\8H2,aOJN-/JRG#QU@_N,c_a<dG
4-=J4PRdEX:V7g/-dE5_]OI2I?Q-&a\F,5G=>FIMF\HQF3@Q0:]5J#;g94e+b-.L
<f;H<f4R.L&NUG).Fg]aCK-+e?WL6Nc9?.T/+-?/)/NSR0b2\&?W1O>aXNCEdSML
(-(cR4IYBR-Y>#g(3>KZ4>^5Q<4Z_e>T+_8B73=aQB3Y>GFFB,?6>[(c#A>5b<X@
PJLf2@_c;L@1D\_K#DZE[><7F40[5cL;15YUc_GDD0eeZ1\=T4_BD<^[d4YDQaV.
(7)[Q6QcXXX<.K+?H/)A=TS@-C;(0@3.a#7c,2gNWFOQX#^-1IMQZN(2>LM1E&C&
8&aYF[PG7K31N(d/O8^KH=#:-c3&QBD8>YLIMJ,ROO\2fd<C+I+PfE_Q/IS24_R;
FIO<bgaD0_E>=D270P(/gK>4EVb,S17W6VZT]A]<AdZ.^)9SN73)X/W5J9&A8HMS
dI)6S/QY:TCF:583PG\VH1,S8<ZR8Z[;^BN:8\T+LR<)EC99Ca?]I,^#2EfKCQM>
a\.8VJXHG@HXa_F#_K)=T-7.NMa+D02@[NV[3P+YR[acT1W[aSG/S]FK#93;R^@R
2+R5=),./@&dB=ERL>4UCUA(Pa,>/U&]LUY,2G3f+5+P@5LB>>L?-?SOKA_U[--1
,gdKG?UIW7FM)>2#1PQOE+QQD4M?T\H5Y)IF2d5+^G3\5KH,:18+ND=Y]^;/])BM
_0F(F+bf-(NYaMa5]DH,RG;CX]EZB\bcM>6fFX#>GJ2/J4_-W9KY:(IR#1aBO>FC
K67)+[4J6^40T;HG+Y97Z<#O)4X0^V>[fMG+PY\?9Ica4.HS.[1K(NgGK382JbPR
G?797EDXg,ZAGgCF,:?W/H,WI+:<Peg_Nd_8FYXR+X;_/ZN34Q#95.=U(Y0(+gW0
89->X@d(T4YQ6<&5VMO;=Gg;QTaN5I,Id9f^X+?8P\4;b9;XLS#Y;ZbQ1>DQ5@)b
>[DDD19/5&+_CJeL1[X]TLQ#d=3P(E@W.X,WL\IUA^Ugfe>be)-_2+gH9?FFQ?+-
W\_d^:OZ6bH#GXb14K4A@37M)40AJW;KWQ:a7K91;I4#5e(M;A<:5@-ZQd<86ZQU
.D[Of>1;<@<JMIG#LMeNL^UfL/,V0K1MUR^61--^IfYCFGHMDed/8UFgUc]T:b7F
P/.WBKBKJ./0VZZB-^;613#;EPfE>LA-<9Lbg0,>.+F8<A+T[DA=_/PPJA)?D0E7
dEd-If5,8);P)a(X(]:5I(E0e?+-<=A7WC/&(PQD_dW)545LF2NKgc7EDOQ+69K[
ISV2#KYV<C66U=V/[Q@&dONJV\N\<@9/Sg_Me=HXR4Q:4V@CL@=VY@Kc^Mc/:N2E
LE,<b?>B66T)V+-cRg<=9JZ;UZ5E86(3Y5OBa)61_@-dUPcK4#5<ITeI^5Z+O1=[
I8]7gX9bQUBD#cF<<^22Y(98f+.A:HU-Z#B75XLT_LJHT&DDO&NTSe9SIUZd<-1X
g->;@R1Lc)_[KE5B8UeP[VW/08Z@S/NIRNbIH^7e53=:5X<OO/-O<1(b@^(G&M+A
FDBRC<J5b@YA?V7((?N8Z06HEfE6]AJJ[A0SNN,G<\@<MK@IZ-HNK(SEQ92HH0aW
([[<J098KD;_Q3-)9bS\T^4Z=^L3QP55HA;/eF_(a^NQ<M@Pa-IA;6+;b;M5BF#Z
OfgR[4@9g1^+@5bSa@OS0(R2aZ^T>B006B1a2-VUfFQ<N;1),9;cE10ZW:DYUgGG
QS:+c6VVfM@_L8dY@=_LAHQ]N6S2+^11W&DM+HVEX_QSIeBE5J9WA]M1V5&G>T[;
:/+LT6L<=^2],I,V(U?((fZW((E2NY#8:94;?6.AEbfLR.-=QX9(8KF3c6Y7I0Ua
BYXP,a??MED:6<GLL26LYR2:FV.>F+S<7TIO70:;^B5BcFfJe]b()_NZd@L\fIMP
,=>,>^_8a19,[?<XWT#6+OVX2-BUAObdT:XgHHU<:(X@McE9@T4)(IgBS@aP6PZY
AT)@B;]SYBVW-KVA(Ib4_BHB<R-<FW,<I+KGKAWYA2a:SQJRaLF#V+&&OcK98#(K
/],NBN0ge&F1+-5d+6Zg(TM?(50Y7D@F[M76EC:e<257.;?4FdO7/bP14A3[+9=U
03;<:6:_\^=Sf(eC@]EVf[Q:OgaLE^#5>;=Y_M4-B?fDW(U2W>8TCYf8[FEZA[1#
NdXeY5/NU4LN3L&41AIW6&0dF<X@(A8cK<FOHA)a_)dDUNU&G[S>-C5,:0GY:9;Z
Q4J;EZa->P<_W^-)LaXfaVIC,9Y-UgcRZMB1Be8SD@(#Z&ffFP((gC[&LeV<g2]1
T28XMAQ,Z[;C[\[G-2=aGOJMJPAQfVYc-Q)ESBc[>UE#,AA,QJ4SFW[H82C@>>_.
CY1DD3]BX2-8A++KHVc#&\&,L/L[>[Ped22WJ_1W;120.8M4E7MBIGIX,)])FgAX
Ygd?.B@1J;97g[:0g\P[Yb6Ad,fC=0;CPg[W[d>)U\)><LZCI+KbfH)9ZFVVWJX3
aS5FZY.b?HGZHeBBR>3?Fg\-C&aUAg6U5WDNE7g+@RSXIGD#YeTC<SXLI?W@+9AX
GPL@&KK>1\4)8;/S]#6R2\aX-EEZg\;7-cT4Y17f3VP:C]T@Ha=FKe1Q4]K8RFTQ
b<N-<=aF96/R=7KF9Y-Q1I55b^L>MM1AXJ4=\G(52<T07WBY@=/=CUJ2+J2^,AEL
E#CFN^_bBGB)&gO8R>6RHU[1J,c9<]eJ^H]C/OBI/6UOAQOGCW\1OHUa)7Zbf^cJ
Cb-fF>aJ)#)[,&3e&U11-@MM5GgV3dIJ8>#Sc)2X.QdW4bXL1K\a00&#][fO#ffa
^f9g#5a?<)@2F54CEgHC3b:C8M,UT>BfX@??b&4+;P7dRD=WQ@3VEEaPgHL#fQ7-
_\NgPH<dY]D:Q?eM2OYB=/da.]X9D1B4a(DP&c/#979f)@8_+H<6G@@PSH4<Y?DT
R#T/(HF/,LJ#ADMP[S&8O?=U?:BG#SU+=fXeXaI)C0G]5/EQJ;)C6-TLXBNW7OZ]
G)X,#BFga^>IVO5VcG1S8A-.UEDA/H@)#)WWNBK4M[NS,CfU@]eSbSJgR+FWE;=E
Q0;&JY1)@C</+:F)TFbMA+;);X2TL/B@JD.cdS-99SV);eJZDgc]NdXAeG>eQ/BA
H8MF-Y.^:D2e>IT\MM9OX+KP+2=5FL9X#2dR@?,d6WaR?:bV]5C4UYR^-UK()VSb
S1VV)-.DLH#DM4-R9AE:Vga/7GCR]&N.:QcIgO>5Q.4e[H/E4O=[53eI[D3LS2d9
KSc&?<=DA&9/cTcUCL-ORGRdQ]:M<,0R6+FFP+Xe?YV0-#&BRKN7R(^+DCgO6R+(
^8C4G-+W,W/N:BJT]1F3<MY(VUH+e)gOVZQI,T[,Kad)FX:[fc+[B:VKg_4JZ[.O
a4D#:/gLa4;JI.:P&MLHg70??Q#IK?<-\FG4.@B/V(K8K:eBJgT/<;J(?.T(-2LY
6g)IfGN0JYUaYJOL&\10_FU7Ba::\Md5=Ae=.]0?O&e>\b/C2gMBC_NGRSbT)OCb
A_,63Ee(42_FWRJUFP?R=CJe4&TZ2EW_=BNOOP,KUaK[+aSXBb.<9_8)aFOXXQ1G
EB1U]W9?6;C[b(P7GMLeM-<D[??b_P5C1f>dO^:O8@L2T8cSNELO2MG=dS8EH,72T$
`endprotected
endmodule