/RAID2/COURSE/2025_Spring/iclab/iclab023/Lab11/05_APR/LEF/SRAM_L1.lef