../00_TESTBED/pseudo_DRAM.sv