`ifdef RTL
    `define CYCLE_TIME 20.0
`endif
`ifdef GATE
    `define CYCLE_TIME 20.0
`endif

module PATTERN #(parameter IP_WIDTH = 7)(
    //Output Port
    IN_Dividend,
	IN_Divisor,
    //Input Port
	OUT_Quotient
);
// ========================================
// Input & Output
// ========================================
output reg [IP_WIDTH*4-1:0] IN_Dividend;
output reg [IP_WIDTH*4-1:0] IN_Divisor;

input [IP_WIDTH*4-1:0] OUT_Quotient;


`protected
<61/\,?<7#Mf#3OVf4XNZS&(SMeAMVDbE+8:6)@#[NW<X@1]/N#8&)d-380\O^[^
L?SXc&<?H4&X;AA-X#IL4.3W061@+Jd=6;))AAO+FJK;KN)#Z]b&b=0C9WW@3BHM
TcY6>.XMM6Y]^=YR_]A.].L&XW<:V[99VCaA7FSb==<7FOZ9#HD^W:MKOHTEV2YF
dU=R/-^<Wf6..,/H>DJ7\3DU2b,/TURgYS^\(1\(d/1A5]T<;I<\]<0@:(6>a@+g
1]]Dd>]X,IPOC9N7>F-Q[GFW]YC>UN[D/./.VbH3aBE@9c9Gb(SBZ18e);76V:#d
0(GRe4OZZ-(9dILN/Oc#EXe2\5Y_c.N71C=79T?Q-&=;74,HE66Y-\(NWKYG5(C6
E5>+OFVS1@)B#S9(@e/A[>II=dQ?CebN3;-JC;)/AH9b)HRcEW)[cHKZ=cZYCQUB
^E3JeU7HWMQA-_?]-#TB<XcVaRdP0U^Q?0;;W[OWf8SM\YN8+66,#3+OP7OSY1OZ
g8XI^OP9Y@24&DW\R-_I(G<XBc>dfY(=6Z/DWY+85CGC\59)Z@G2/#>Ef(QN/V>,
gSQX<SbY#E([8<MOeN<+5_(@VHCPfd(LBDEgeX&^)/6f?G+c@@[[#CNJD6B+8ZN7
bP)(E7=D((N2VV(Y5Dc:eC\&>KEE0cb:2g0QJ#HA<P&&QCC/L3RQ2F9P-+f5.XeI
J@,Z:.G^?V7)JP=.,W7Z:XVVO\AB)6Q[H<3CZ[e_KSI+aMbZ3S<>ENGCK#QHC18A
F@V2=S>b/AYdHFAZB+=[8fbKg&dZ7Ie;LF5;E)Te(5=G1MW]C?68+^1IIaU;<KPb
(UPH(16I.bLDQWU.3(0C@OF(7CE0Z/P/6\TOZ[N:,b5g8[eTMA4>5SLP/>+),c1^
gER4?V(:)JQ_Ma8LgZ[WQ0#A7WR9C-DZ]e.VLA,YPeb<XgS4C/aU/:4bA>6I#@=>
dAgS74@URd[dYcXR5McZM+&_=WE&SB5P:)T(];&0(:[9()CKHfCaREH@BXIYO\23
bP4=dS]C0RVG^Pa?Xfb;;O)?76?P1[G0TWgBS9,S=OK43[OG1&0=f&<aV>RV@M.7
_ASb/cZC>FZdM_#=N>;SYSeCG]9Z;MPX+DA0=ICJI9Z;T>ND(E7^PK02?^&]VGVY
A7@.aA&dd;RE<G+B#ILSHe)HOEZH:A_eA<Q^<b)?NNdJATK?R6>-O,gF\Y-4=(E<
+N.R[c@c<NM.C9F](a^SS/a:PIM@NE#]M#bBGb:@4Z-D&G,]0:SHKC:+5RWTEK_D
I??c5d6=\#)Ge<D3bY5X0N\KG+6?_B-))g,N)MeN0WBJPX[=I6ON2;#</_W._4[9
\8@J_WVD24BJD8H/)R+N5#R7b(FO+F5_]3]^@B_c/-9^B<)+^FP5\-FHf9IgG+1Z
N5ePbNS2^+S&]c46AT=.dFHY#-_R9MV_E1W&IJ4U\8>#C<#R(Y>g.+I_I-DZ.aFA
G<aZCOb6PBLFBGb6:KKfc))^B+HAMUA5g)_K]2CVf\W]5A5^21LBKAWCXZO[P9;E
X\aNf4@GME;^^D\a)^[fH0,bOV(]\BM;206)7]ZHSI0K)O&KPg4c8=@^,GFbB/RR
>K2+:V;><:AT5<^^H7FBOW,VeHFMD3Z\9bCEB2J+:G/8?)3W>B>RJbf8g+)81G+0
,DGG-B&[K6>d#b:OHM/#+(27.(URQ1Ce^<^bYM1G#X?e+(Cd=7#0@fKPeVJ;A.1E
A<_<^738CSMN=+[9;MbGgf7^GG5TB/.Q6W[V6\PMXZ&VAAKE,-13OX)HUaS[=FZI
S6B-#T#b8EYUGCY8]bIB+\2EZ-BSJ(YAAR)#)X(W+X]fO^5B&IA<>+ITP0U1JO0L
f;T1cb+UeY>T.VaV,\#.b.]3S[A,gWX9@R=#Rb]ZT4OC;]YL@71U#b)\R9^YecXd
)7J<.T&K(^S;3gI-bQNZ,?2NY-.T:6M[A:]25M@RA)B,82-:P4^Pd&_,e96&0FZT
Xf,0ZD)aI\V7]\WX&9F)MSV9b/d=6@[&9#,T3@SSF>dU(?1,R93fXH^f5W(4>Eb]
bOTF<<&D&UaD?dBKCMa2C4bd=;ZSaA.QgV?D@Q^7CgEPC,6fQ,7]T&EO0;)(@PVY
J?Q;MWgWfMdb=[N/3#202HQ76Y.Le+4Y19BPL]9XM^#A,S,TdF=^Q>K\T-DPNX[A
X?UYMRS]c158(BUGGO@FG_T.Z]eV.&Y#UN&c:@(YV^5b51>+IH:7CE#X47Kg_/3>
#EB](,V7#P,Q6>d70]JXGIYVS)V#Ld0@@:493:fTW=J4Q;T,8I]2CQDU@V2XG/SO
>OII-A:D^]c.e66V5+2IDOe=Z)HHE2L5HJ.#YG?T?S([cH,ASWDG=7L)94;TNQdC
[)6;fFN@\X0CN)XQHC+>-EcaVZ.0Yaab0LN?<8)(WU.?=/@;c^PL\Rfd/2Ng-e+1
234f]+U3O<>\UQGDJ&@0dcL]+(H-N^>g//5DLRY5=g:aUgCbe]).+6SDeaUbZ?I=
8K)QASeNB1a5+]935U3,C3.2]S0ABA,\\b>U=V6=+IFYdW<-,PR/1De3+?H@&9P<
YV/ZXbIVRA3MT&5,e3gFH#,)-Te7#KZEW95#P0R\,+-TA,>Ug#)<-K[QfR@_c&<2
R?()d(K_MF0dN)LE&2\_YQH(XH7EI@CF6>EH?/:ZS_N5K&^g#/R4>1OfC3MS9QA/
N&(.SgGgMfNbZN>C9S]I&#g646HgE/VJ?F?Yc-+=EC;cA-5N<40,O@=+9)+0KA=[
H)D:O:>8W?IS<Mf97LJD>BNeg;Z@6WS>f\V11]NR+UXe.0Q=Y(-;+fc=&O3#9?3H
\S&c.E95.bP&gbea0(8aVP=MKF<Tg1Y^B3GFM)eV5GOS(F^KH-e+AK_H=N60&L(9
8d+_0M2Y::Wg6?OI=e-4W(EH<M)/JH&)N2,:A[\,;C2T<fP7cV><J@^T=<g\,W[-
ULG7+Q3/F0LNb6PHeD)XHRQ]E0-C=c8F_1-b.(.94b_#TgFS).YL)eM^D12;+gC/
,]KF5?C<7UJ9=UbE6=:.&9c#T:.;;eTQM>AMLC7Y^OUVC4:^/(:&MV-/SW)-&>&Q
OWAB8Q&._=Pd5g(8G7M)X89YbU[QF[WR3&P^;>.7M@Zd]T)>?@KMY0W_C(VEL)8/
FW?N,#d,XZFVE-^4>NcEE0;dJE&X84WJ:\>A.N>DM=@d[?B;gB\(G)^c7G/FG[E:
+QCK0AA;1IKLGE7&Oad?UECa/\gJA1T7Q1>eDRfJ7U0R\>+0/A(44N.Ie_NI(U3W
&W8Dg5438BG\MP/C,H??g:KIc,B9/3e2Q>:WDeUN&:(#N]MC8U<5/5/VTGg=&RM-
O]Q/)&FQKRTfA2DSZFE3GVKCI,:Ob@SDIW9AH0dc6XNI/2O/]@E+,8fUZ4ZG>X_.
1DRVW&8BdBDDP#5-2XVVEgXbY0_6-PD_W1OX]g(+QVP)7a+1g<6A(d@:_EY)=.;>
S3V?1adcc&7#]gZ4UcMF=gcK58b9Q<P&(LX2-C,EO[5.^a[Me?GfZZV)X,9L2,47
R]5I#V>5H84EY.RTCL:TDPJCdRH3-S6g#<@MQ30Yf9#G4,^LPM\G^Z9PCdIB@V&\
-gF0ZXNKW3^RC;fSODQ0980f(:b/Gg7NL8>](4U2Nf_N_P:A;?6ZcS9=5c7;c.>K
>69@OgCEBIUK^(I/CYgMZBZOT^4LBIe#8=aI^]CXE(2AYU=)7;fYW9?/JGXOf-aF
W2G3&d@I6?)4@@ZZU]6b;9Z([;+dG5PTKLY#MTCTU+&?1d\F9OX>ASdE<39=:K+d
+HRXG8cSe/b#6#(#\H)Le\J>\D)M8GNRQDB1?gXX<->=[<?-+L0QHeA2DaDd8175
IN1,2Y/WG1T&.7f,4]#^\@TgT?UK=B\2VF]BOU)W@a/J>9QBK+8g:_3ONR+0#C0<
7=[2A@1JdH/>K@(+@(RH=<LOV<_Va\C@g3.MOgQdB(e8^D<V@PZdUg03?H>2\C)I
#216M;8,d?,FBH[;YN]<_#B+&0e^RH_dA&(HbE>O=Y6B]gBcRbC,C>-B9FEK_SW7
28B,b8>9Y]HWOKT31aEgTAW6QMO>A,4<TF.f]b,LT4:QeYGN(AW9II@&POBf,-FN
C=M;NGeaJ.g4JN7F/]5G(]_,HVZ;72.@1e.W(@&RY2^fH\KY^N47M9RBd:Nc>&)#
#N0&Aa[LL6(04M>/]5IZ?-c&IGRE^LV:Cg2#0b9#AI+Z]EC0Dd_K0>@/583KB)T@
H(6N>K^&@9@HK)9Q@7Td=D@Xf,ZD8,Q]_DC^)9d+5R#]SWNcG[L)USf7QKOIe52J
+?aK;K?&UO.]Y7USN3-OdTfM8THdD^XCS.g8&]5_<PD_5M:F&DIRbO-[ZXeJHGUT
CQN07V#TU2/cG/:6dgg)/A7&:9MHH^U5)XH6GJS4fU#9F.EB+MZ<\9N..fdSV&]c
-=X@(>;5[]6fFDU517c435&G#?,2;G+IN@R/LK3:dSUXaN;>B]FU1W9H:XdeF)79
gf58E[^DWQ?MOG@YXd\8E>=ZOWbHZ<6A?CTdc:Qa(CO1GHF(==BFVGZ-fGP4T:U[
)fZTcEWD@]B4f1R7?)PYX=9f\b.6:[fGYY5KTVN\eWe1:.UV0:Z.3a]6I,Q@+-Ub
NSgH0PJI=.TBDIT\+LPAacI+Cg=.E[G,D3cZ0IN^.?6BP=A?UB1=J;5>fd7AU8_E
YG.eN,M4V:PYS:H#HAYNc[)f6VQVNJ\d0-?eF>BSPSUMaO+,3?9I[6bSN_I?IeG>
LUQ/TY(?E(cZ3_AH\2S>9RaLN2V/fD91K;4D4]G-LO)B/_\>IBJZOEUT.?Z,4)?X
.D^eZUVeC_c,HU(:@?MFX-S&f1bIc#SN+1PG6M)R&/_0DY+1>WABJ(9D6415P:cI
&;)0:^Y9cIV?Bd8Q]<a2d,,(J/)4H:8>W2-X>J/4:X@:?g_,[R<J4,A/VU-GT().
X90K-@1@\\W7EZGT31Z07XW58\@;SJR4a7K2@AfNDd\/&.f.dA[XV_KB+(RfOUYZ
9T^MB=8,bfQ-L9@(6a2X&[cg-(11Z?G/Y^<O5<aCH#&GE5MgJ-fK]b,]&<TTa4D?
>N?cY3,5P23Y_-3<BN7eBP+Vb/M)QO#QQ2A5&\WOK(cG(+,)D(8H08N3Z[:;+8=1
N/CL<Y\/GB(Hg&E8C=;8W4>0IAB^:PIVdY)UQ;SO2/7;-geLG^#WbJ=/gA@6>\?c
[\;\-Q&MXCE6QaV@==AF@#BQ.#))9/ZSF<IF:/MK]A\VFIBF,dK.fNHT^6NFBDJ?
UQRdOF2XPN3D1(RffXb.c2#]P?_OR028GV7(cEF(C8@APgL8Tf-M9Yb+K_C65)J3
UeKDSJdc[@:UKWVPe(?\NG)=KW7?6&#G2aH^J9)E50Y+WPZHW@?300RWX,8]?c.V
XMT;0;=g&<ER3LYL&M-3L\HgQCR>8P::N\K^-LIGQ5K.##d0D4V,W;a#>Y6HBR3/
X#8IN_b2SggR2Md:=HCEK[6gXY0J+;8YY?3#I[L<M;I@=)#^cZHVY/BBT:<HW=EY
CWeT0)4LXK^>ReSQ=VC.QN#04Je^4cVX>gM=)QJG9B,]\E4GPgY0^VT=)Z72b^.#
g6^,H1(NRdK(XOcPgNZU<e>5+LZV1AT(-=14a[W-68=<0=BZ,b&g9^7-K_8JD[-g
45492Y-7?K[bWDc41+K\UP&@c@;N)M@Ta<J,XcV1J_b0ZER^Nf6c+/;L^_JE0b0W
3\+-I<FR_&)KPFV0MI0E#\WcQ]IA0E\]?$
`endprotected
endmodule