../00_TESTBED/Usertype.sv