../00_TESTBED/Usertype_PKG.sv