../00_TESTBED/PATTERN.sv