../00_TESTBED/CHECKER.sv